use WORK.ALL;

library IEEE;
use IEEE.STD_LOGIC_1164.ALL;
use ieee.numeric_std.all;
use Std.TextIO.all;
use work.debugtools.all;

ENTITY ram8x32k IS
  PORT (
    clka : IN STD_LOGIC;
    ena : IN STD_LOGIC;
    wea : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addra : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    dina : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    douta : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    clkb : IN STD_LOGIC;
    web : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    addrb : IN STD_LOGIC_VECTOR(14 DOWNTO 0);
    dinb : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    doutb : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
END ram8x32k;

architecture behavioural of ram8x32k is

  type ram_t is array (0 to 32767) of std_logic_vector(7 downto 0);
  shared variable ram : ram_t := (x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"20",x"01",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"4D",x"36",x"35",x"55",x"43",x"4F",x"4E",x"46",x"49",x"47",x"55",x"52",x"45",x"20",x"4D",x"45",x"47",x"41",x"36",x"35",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"DA",x"1A",x"0D",x"08",x"50",x"08",x"56",x"23",x"01",x"08",x"0B",x"08",x"37",x"01",x"9E",x"32",x"30",x"36",x"31",x"00",x"00",x"00",x"BA",x"BD",x"DC",x"21",x"9D",x"FC",x"00",x"CA",x"D0",x"F7",x"A0",x"35",x"4C",x"8E",x"21",x"3C",x"82",x"06",x"B1",x"34",x"09",x"C9",x"6F",x"0B",x"34",x"0C",x"59",x"A9",x"AC",x"05",x"4A",x"4A",x"03",x"28",x"A7",x"FA",x"91",x"0E",x"01",x"0F",x"04",x"00",x"7E",x"8E",x"81",x"7B",x"0B",x"60",x"B0",x"60",x"6E",x"B7",x"CD",x"F6",x"DA",x"03",x"0F",x"02",x"02",x"3D",x"E1",x"F3",x"2F",x"E6",x"76",x"DB",x"6C",x"AF",x"3D",x"0C",x"60",x"0A",x"07",x"AD",x"0D",x"15",x"0E",x"28",x"BE",x"03",x"83",x"27",x"85",x"54",x"70",x"19",x"D7",x"4C",x"5C",x"F7",x"98",x"AC",x"EE",x"B1",x"6A",x"FD",x"37",x"3B",x"6B",x"6D",x"59",x"E2",x"58",x"00",x"26",x"80",x"2C",x"A1",x"2F",x"86",x"66",x"13",x"4F",x"B9",x"DE",x"4E",x"85",x"31",x"2E",x"30",x"E8",x"33",x"01",x"09",x"E4",x"84",x"9F",x"83",x"31",x"62",x"44",x"8A",x"A2",x"06",x"33",x"2D",x"90",x"CB",x"1A",x"A1",x"05",x"89",x"2F",x"46",x"A6",x"DC",x"D6",x"00",x"E4",x"42",x"27",x"BA",x"45",x"86",x"63",x"09",x"00",x"EE",x"CE",x"00",x"2A",x"12",x"0F",x"27",x"0A",x"B4",x"D1",x"BA",x"5B",x"F1",x"81",x"9B",x"02",x"17",x"A3",x"ED",x"72",x"1F",x"24",x"78",x"8F",x"6C",x"36",x"E7",x"50",x"3F",x"1D",x"61",x"27",x"06",x"56",x"CF",x"95",x"1B",x"F3",x"CD",x"C4",x"5A",x"30",x"DE",x"35",x"22",x"06",x"92",x"E5",x"6E",x"20",x"67",x"C1",x"30",x"3F",x"19",x"C1",x"95",x"CC",x"84",x"A5",x"B9",x"1D",x"3F",x"1C",x"70",x"B8",x"6B",x"05",x"2D",x"B7",x"21",x"89",x"E5",x"EA",x"6C",x"78",x"00",x"31",x"F7",x"6E",x"AE",x"26",x"77",x"2E",x"09",x"3C",x"1D",x"3F",x"49",x"A1",x"DA",x"5D",x"6A",x"7B",x"3B",x"92",x"E9",x"64",x"CE",x"C4",x"1C",x"41",x"67",x"D7",x"1E",x"F5",x"24",x"5B",x"40",x"CB",x"6C",x"86",x"DE",x"21",x"26",x"C6",x"FC",x"6E",x"E4",x"CC",x"09",x"6E",x"92",x"06",x"47",x"54",x"06",x"9D",x"6B",x"E3",x"CF",x"8C",x"D8",x"62",x"6A",x"30",x"19",x"B3",x"31",x"86",x"33",x"B4",x"0A",x"A6",x"9D",x"10",x"A9",x"66",x"9D",x"2F",x"72",x"16",x"FA",x"50",x"2E",x"A9",x"25",x"65",x"97",x"BA",x"29",x"75",x"C8",x"48",x"32",x"39",x"09",x"55",x"B9",x"77",x"68",x"A2",x"DE",x"1C",x"E3",x"84",x"4F",x"8E",x"49",x"32",x"2F",x"66",x"34",x"F4",x"4F",x"51",x"30",x"C3",x"62",x"94",x"35",x"77",x"2D",x"6A",x"DA",x"75",x"68",x"26",x"18",x"65",x"CA",x"F0",x"F7",x"72",x"94",x"6E",x"70",x"2F",x"A7",x"6B",x"77",x"A9",x"08",x"2C",x"DF",x"E2",x"F1",x"95",x"F5",x"21",x"48",x"45",x"6C",x"1B",x"D0",x"B4",x"15",x"E8",x"27",x"CD",x"8E",x"91",x"73",x"F1",x"A4",x"63",x"75",x"91",x"0C",x"38",x"73",x"37",x"1D",x"02",x"2E",x"8A",x"23",x"BF",x"19",x"D3",x"84",x"79",x"BF",x"D6",x"19",x"99",x"56",x"8C",x"B5",x"8C",x"76",x"98",x"33",x"6C",x"4A",x"56",x"17",x"F2",x"62",x"59",x"2C",x"A5",x"32",x"05",x"EC",x"E2",x"BB",x"E2",x"88",x"2E",x"24",x"66",x"29",x"AE",x"4D",x"70",x"86",x"28",x"F4",x"46",x"CC",x"81",x"70",x"B0",x"FD",x"3A",x"82",x"15",x"79",x"2E",x"E7",x"54",x"57",x"21",x"65",x"8B",x"22",x"35",x"42",x"A4",x"48",x"FB",x"46",x"98",x"6B",x"D8",x"0E",x"EA",x"85",x"53",x"32",x"A8",x"53",x"61",x"78",x"77",x"B5",x"86",x"6E",x"54",x"64",x"4B",x"6E",x"2C",x"54",x"B9",x"AA",x"07",x"21",x"63",x"53",x"17",x"A8",x"37",x"BA",x"00",x"8B",x"4F",x"CC",x"4C",x"D2",x"0D",x"EC",x"0A",x"12",x"7D",x"33",x"26",x"5A",x"7C",x"AD",x"89",x"B3",x"AD",x"16",x"C5",x"64",x"EA",x"0B",x"2C",x"E8",x"C0",x"0C",x"00",x"22",x"1E",x"E3",x"A0",x"48",x"66",x"B9",x"64",x"75",x"6B",x"A0",x"90",x"15",x"50",x"8D",x"21",x"57",x"67",x"1A",x"9C",x"21",x"24",x"68",x"99",x"24",x"D4",x"77",x"59",x"B2",x"CE",x"D1",x"08",x"67",x"98",x"BE",x"4B",x"B7",x"D3",x"68",x"D6",x"D3",x"10",x"C1",x"51",x"B8",x"21",x"67",x"28",x"DC",x"BF",x"13",x"8D",x"88",x"F0",x"04",x"27",x"47",x"6D",x"DE",x"74",x"EC",x"25",x"68",x"04",x"33",x"17",x"B7",x"62",x"71",x"75",x"69",x"9F",x"2C",x"29",x"66",x"97",x"1D",x"6B",x"1D",x"2B",x"7A",x"2E",x"1F",x"70",x"38",x"B5",x"61",x"76",x"36",x"BC",x"9D",x"CD",x"D5",x"C6",x"79",x"A9",x"A0",x"72",x"DA",x"4D",x"E7",x"7A",x"75",x"56",x"7E",x"46",x"9C",x"1E",x"BA",x"E6",x"C8",x"AC",x"D0",x"12",x"E1",x"88",x"79",x"75",x"14",x"18",x"A4",x"C8",x"0A",x"3F",x"65",x"2E",x"D6",x"C3",x"52",x"1E",x"75",x"9A",x"EB",x"21",x"C3",x"AB",x"CB",x"D6",x"2C",x"1A",x"E3",x"0C",x"03",x"3A",x"C3",x"97",x"FF",x"80",x"00",x"02",x"44",x"01",x"B3",x"31",x"C1",x"04",x"04",x"60",x"31",x"83",x"01",x"1E",x"80",x"A9",x"02",x"16",x"3C",x"75",x"90",x"25",x"50",x"75",x"06",x"6E",x"CC",x"E7",x"49",x"26",x"15",x"B7",x"40",x"BC",x"02",x"47",x"33",x"35",x"34",x"A8",x"3B",x"A6",x"00",x"AB",x"05",x"AD",x"77",x"21",x"6A",x"6F",x"79",x"FF",x"F4",x"81",x"78",x"90",x"32",x"11",x"5A",x"25",x"4E",x"61",x"5B",x"8E",x"75",x"4A",x"D3",x"77",x"38",x"8D",x"43",x"25",x"D6",x"0C",x"58",x"2E",x"E4",x"8E",x"35",x"E2",x"9B",x"21",x"0A",x"09",x"9D",x"27",x"8A",x"45",x"BF",x"00",x"67",x"A1",x"FC",x"F0",x"6D",x"B8",x"74",x"16",x"E6",x"64",x"02",x"68",x"14",x"D5",x"DA",x"E1",x"A8",x"57",x"33",x"70",x"F3",x"01",x"6E",x"D3",x"61",x"41",x"F6",x"B6",x"CC",x"5D",x"6F",x"04",x"6D",x"2D",x"6C",x"40",x"79",x"29",x"3A",x"1E",x"4F",x"01",x"15",x"D8",x"45",x"31",x"C9",x"25",x"BC",x"46",x"1B",x"1E",x"AE",x"03",x"6C",x"FA",x"59",x"11",x"A9",x"1A",x"63",x"24",x"E5",x"10",x"1D",x"11",x"33",x"2E",x"35",x"22",x"7C",x"5B",x"07",x"EB",x"70",x"79",x"B5",x"58",x"30",x"84",x"41",x"00",x"8B",x"7B",x"DE",x"1D",x"A4",x"1D",x"06",x"3A",x"01",x"0B",x"E4",x"04",x"00",x"08",x"ED",x"17",x"75",x"6B",x"E4",x"94",x"12",x"CA",x"47",x"58",x"6F",x"9A",x"6E",x"EE",x"9D",x"68",x"95",x"EE",x"DC",x"80",x"46",x"D0",x"EE",x"56",x"12",x"64",x"95",x"1F",x"3D",x"56",x"63",x"AD",x"65",x"76",x"25",x"E1",x"2C",x"49",x"13",x"BC",x"88",x"9A",x"72",x"6F",x"6D",x"7B",x"3C",x"D0",x"39",x"A7",x"2A",x"35",x"32",x"D4",x"33",x"29",x"05",x"66",x"30",x"31",x"38",x"62",x"FF",x"0F",x"D5",x"6E",x"10",x"6C",x"B3",x"17",x"7A",x"20",x"6D",x"6E",x"23",x"6C",x"75",x"81",x"70",x"36",x"79",x"D5",x"07",x"DA",x"96",x"73",x"D6",x"40",x"06",x"A4",x"61",x"B9",x"62",x"6C",x"BF",x"50",x"56",x"0E",x"19",x"7F",x"D5",x"02",x"A6",x"D8",x"0B",x"6E",x"8D",x"95",x"AF",x"3B",x"3A",x"13",x"DC",x"70",x"97",x"22",x"AD",x"2E",x"05",x"35",x"37",x"A7",x"14",x"6E",x"6D",x"9A",x"87",x"60",x"36",x"8B",x"68",x"7A",x"3A",x"71",x"37",x"32",x"8F",x"2A",x"34",x"A6",x"75",x"8A",x"0D",x"00",x"02",x"0E",x"FB",x"9A",x"67",x"65",x"0D",x"5E",x"20",x"3B",x"5B",x"CB",x"E7",x"3A",x"15",x"5E",x"74",x"AC",x"98",x"8A",x"D5",x"6A",x"C1",x"14",x"97",x"13",x"64",x"61",x"08",x"CF",x"9D",x"6C",x"D2",x"C3",x"28",x"B6",x"2B",x"43",x"29",x"C6",x"21",x"6A",x"73",x"0E",x"63",x"72",x"5F",x"77",x"65",x"6D",x"37",x"78",x"57",x"E3",x"C0",x"71",x"82",x"0F",x"AF",x"40",x"0D",x"32",x"3A",x"C1",x"47",x"70",x"D9",x"EC",x"3A",x"06",x"76",x"12",x"04",x"6D",x"4E",x"6D",x"CF",x"22",x"32",x"0F",x"73",x"EE",x"D5",x"B8",x"67",x"36",x"84",x"9A",x"61",x"74",x"6D",x"C2",x"6E",x"3A",x"5D",x"36",x"C5",x"31",x"04",x"0E",x"35",x"38",x"30",x"3D",x"2B",x"0F",x"9F",x"77",x"68",x"70",x"53",x"D4",x"A8",x"A3",x"5B",x"0A",x"63",x"B6",x"68",x"6F",x"DD",x"54",x"6C",x"63",x"02",x"6E",x"EE",x"97",x"79",x"28",x"CA",x"E1",x"01",x"10",x"64",x"4C",x"67",x"EB",x"5C",x"B0",x"6D",x"70",x"6C",x"3D",x"94",x"69",x"65",x"72",x"3A",x"6C",x"23",x"66",x"02",x"D0",x"9D",x"4E",x"94",x"03",x"00",x"80",x"0E",x"64",x"FA",x"3A",x"6C",x"67",x"E2",x"92",x"73",x"8A",x"3A",x"E8",x"64",x"1D",x"49",x"70",x"77",x"AF",x"90",x"03",x"86",x"7D",x"10",x"50",x"06",x"FE",x"0C",x"6D",x"75",x"E0",x"48",x"0E",x"64",x"28",x"50",x"73",x"3A",x"06",x"08",x"00",x"9D",x"83",x"13",x"AA",x"92",x"77",x"11",x"CF",x"68",x"75",x"D6",x"BF",x"71",x"85",x"8A",x"18",x"28",x"73",x"EC",x"21",x"83",x"3B",x"63",x"96",x"72",x"B6",x"79",x"99",x"0A",x"10",x"1D",x"7E",x"12",x"46",x"72",x"65",x"E3",x"B3",x"29",x"24",x"74",x"54",x"20",x"54",x"84",x"62",x"6F",x"5A",x"72",x"E9",x"69",x"6E",x"67",x"EB",x"10",x"19",x"4F",x"43",x"76",x"A7",x"D0",x"CC",x"58",x"4D",x"66",x"75",x"A7",x"6C",x"97",x"73",x"8E",x"48",x"64",x"20",x"FB",x"78",x"69",x"74",x"00",x"F5",x"38",x"06",x"44",x"61",x"6E",x"D1",x"63",x"65",x"6C",x"87",x"19",x"00",x"B6",x"3F",x"20",x"0D",x"30",x"11",x"0D",x"20",x"40",x"10",x"02",x"6F",x"6B",x"F8",x"37",x"A3",x"11",x"56",x"C1",x"8F",x"F9",x"46",x"14",x"8D",x"18",x"D0",x"F5",x"78",x"20",x"C1",x"31",x"5F",x"10",x"F7",x"6B",x"71",x"F8",x"AD",x"FD",x"75",x"F9",x"68",x"0F",x"FA",x"AD",x"54",x"29",x"AD",x"29",x"6D",x"5E",x"40",x"EE",x"AD",x"F8",x"02",x"90",x"05",x"5C",x"5F",x"FC",x"BE",x"DB",x"12",x"D5",x"47",x"63",x"40",x"E2",x"C9",x"67",x"FD",x"8D",x"3B",x"BC",x"33",x"4D",x"0B",x"47",x"0A",x"5A",x"CC",x"D0",x"04",x"18",x"97",x"82",x"4B",x"B0",x"0A",x"B1",x"AB",x"56",x"BC",x"42",x"38",x"3F",x"58",x"2B",x"03",x"1F",x"74",x"7B",x"19",x"7F",x"58",x"78",x"70",x"47",x"F0",x"03",x"EB",x"CA",x"B5",x"D0",x"59",x"4E",x"02",x"63",x"49",x"BE",x"1F",x"95",x"42",x"F0",x"1A",x"AD",x"5C",x"3B",x"FB",x"7B",x"20",x"5D",x"52",x"8A",x"66",x"94",x"86",x"D0",x"59",x"A8",x"71",x"B2",x"22",x"9B",x"57",x"32",x"35",x"89",x"3D",x"23",x"79",x"29",x"E4",x"34",x"BA",x"D1",x"9F",x"2F",x"F9",x"C9",x"F8",x"D0",x"0E",x"FB",x"35",x"13",x"D4",x"14",x"77",x"82",x"42",x"A4",x"D9",x"66",x"6B",x"85",x"91",x"8C",x"13",x"25",x"64",x"B3",x"1D",x"D4",x"F3",x"39",x"98",x"23",x"9D",x"1A",x"46",x"5B",x"F1",x"A7",x"CE",x"F4",x"E3",x"B4",x"2C",x"F2",x"8C",x"60",x"C7",x"24",x"39",x"42",x"F7",x"5C",x"FA",x"05",x"2A",x"0F",x"41",x"1F",x"1D",x"1D",x"8A",x"BD",x"CA",x"C7",x"9E",x"A7",x"48",x"AD",x"52",x"2A",x"A5",x"48",x"5D",x"53",x"51",x"AE",x"94",x"65",x"1F",x"BC",x"F5",x"A7",x"46",x"D8",x"7A",x"1C",x"1A",x"3E",x"E1",x"22",x"7E",x"68",x"DC",x"42",x"EB",x"D4",x"06",x"B2",x"4E",x"16",x"46",x"9E",x"4C",x"C4",x"11",x"20",x"F7",x"CD",x"12",x"55",x"D7",x"FB",x"2B",x"95",x"26",x"F6",x"EE",x"5D",x"DA",x"BA",x"03",x"27",x"55",x"31",x"55",x"56",x"A5",x"F3",x"3A",x"57",x"0D",x"8D",x"62",x"01",x"6C",x"43",x"09",x"B0",x"16",x"44",x"50",x"08",x"C1",x"2B",x"91",x"30",x"EB",x"A2",x"DB",x"03",x"7F",x"32",x"00",x"09",x"01",x"A9",x"EE",x"06",x"9D",x"BB",x"53",x"2F",x"0B",x"41",x"6C",x"F3",x"FF",x"EB",x"21",x"4C",x"34",x"13",x"DB",x"E7",x"B0",x"60",x"AE",x"DC",x"67",x"05",x"7A",x"57",x"BC",x"8E",x"58",x"38",x"8A",x"29",x"D0",x"30",x"30",x"96",x"59",x"F7",x"31",x"5A",x"DE",x"32",x"7B",x"5B",x"33",x"EF",x"5C",x"34",x"BD",x"5D",x"77",x"BD",x"35",x"7A",x"5E",x"58",x"51",x"5A",x"1D",x"A6",x"AB",x"59",x"08",x"F3",x"21",x"D0",x"74",x"03",x"C2",x"1E",x"C3",x"8D",x"16",x"00",x"6B",x"A0",x"CC",x"C0",x"BB",x"63",x"4F",x"B9",x"4B",x"99",x"DA",x"47",x"88",x"0B",x"16",x"78",x"11",x"09",x"6A",x"DE",x"78",x"EF",x"04",x"2D",x"20",x"A3",x"C6",x"13",x"D3",x"39",x"86",x"5C",x"A5",x"42",x"4E",x"EA",x"A9",x"81",x"27",x"FE",x"04",x"F2",x"A1",x"11",x"BA",x"12",x"7B",x"78",x"C3",x"DE",x"FA",x"BD",x"C8",x"DF",x"BA",x"E8",x"93",x"D0",x"F1",x"9B",x"BB",x"1F",x"60",x"AD",x"84",x"0D",x"97",x"D4",x"B5",x"7B",x"5A",x"AA",x"55",x"58",x"6B",x"49",x"C1",x"EF",x"F7",x"B5",x"AB",x"00",x"94",x"B2",x"6B",x"B5",x"A2",x"DA",x"AD",x"DF",x"72",x"FA",x"29",x"32",x"80",x"B3",x"73",x"5A",x"41",x"F5",x"26",x"17",x"06",x"35",x"F4",x"25",x"17",x"80",x"8D",x"0F",x"C0",x"D2",x"0F",x"5F",x"20",x"0E",x"14",x"0E",x"BD",x"07",x"B3",x"08",x"F2",x"BB",x"AA",x"B3",x"08",x"F1",x"BB",x"2C",x"B4",x"CC",x"32",x"A2",x"F0",x"AB",x"4A",x"8B",x"B0",x"F3",x"AB",x"52",x"8B",x"B0",x"F4",x"AB",x"5A",x"8B",x"C1",x"B0",x"8D",x"F5",x"C3",x"7F",x"9D",x"14",x"E1",x"1D",x"57",x"20",x"93",x"23",x"5F",x"C1",x"9D",x"82",x"5E",x"07",x"E7",x"25",x"61",x"B8",x"62",x"60",x"61",x"1B",x"88",x"C9",x"C4",x"C4",x"19",x"A8",x"B9",x"84",x"C5",x"8E",x"F4",x"22",x"DE",x"FD",x"CA",x"D0",x"F8",x"FD",x"23",x"83",x"93",x"0B",x"8F",x"27",x"53",x"F7",x"A9",x"0A",x"57",x"A2",x"D0",x"05",x"CD",x"ED",x"70",x"F0",x"26",x"9B",x"10",x"70",x"23",x"06",x"54",x"F8",x"82",x"84",x"4C",x"B0",x"8D",x"F9",x"73",x"8A",x"FA",x"A9",x"80",x"C8",x"AD",x"F6",x"F4",x"06",x"9E",x"DE",x"22",x"E9",x"CA",x"C4",x"5F",x"48",x"8C",x"B5",x"2F",x"2B",x"61",x"47",x"C3",x"60",x"1B",x"20",x"CB",x"05",x"15",x"AF",x"A3",x"00",x"E5",x"60",x"7A",x"5F",x"3C",x"5E",x"1E",x"3C",x"60",x"8F",x"5F",x"47",x"21",x"5E",x"A3",x"6D",x"AD",x"4D",x"A7",x"4D",x"AD",x"AA",x"A5",x"17",x"AD",x"A9",x"4E",x"C6",x"AB",x"53",x"58",x"61",x"EF",x"59",x"62",x"BD",x"78",x"53",x"F9",x"8D",x"63",x"0D",x"1C",x"BF",x"A2",x"71",x"52",x"7D",x"4D",x"DE",x"D6",x"88",x"7E",x"FA",x"4A",x"6A",x"F5",x"90",x"F5",x"B3",x"B6",x"12",x"ED",x"89",x"27",x"DB",x"59",x"A2",x"49",x"AA",x"BB",x"22",x"AD",x"49",x"C5",x"76",x"35",x"06",x"23",x"94",x"4C",x"F1",x"15",x"A5",x"F3",x"7F",x"8C",x"D6",x"DE",x"BE",x"7F",x"28",x"BA",x"55",x"2D",x"07",x"24",x"FF",x"CD",x"00",x"C0",x"DE",x"EC",x"7B",x"E6",x"A2",x"27",x"BD",x"63",x"F9",x"5C",x"D0",x"3D",x"9D",x"C0",x"07",x"CA",x"5E",x"F2",x"68",x"7E",x"C5",x"B9",x"FE",x"F0",x"06",x"FB",x"4C",x"1C",x"16",x"8D",x"6F",x"AB",x"E6",x"43",x"A9",x"0F",x"98",x"35",x"08",x"EF",x"03",x"B7",x"85",x"57",x"E3",x"8A",x"C2",x"7B",x"00",x"DA",x"C2",x"7B",x"80",x"AC",x"11",x"DE",x"03",x"E8",x"24",x"BC",x"22",x"E9",x"80",x"52",x"78",x"19",x"FD",x"A0",x"14",x"5E",x"EB",x"89",x"4A",x"01",x"37",x"0C",x"6F",x"03",x"E9",x"0D",x"CB",x"77",x"10",x"20",x"DE",x"3D",x"DE",x"ED",x"A9",x"21",x"2B",x"6C",x"16",x"AC",x"D5",x"35",x"FA",x"1E",x"00",x"ED",x"00",x"F4",x"65",x"16",x"65",x"40",x"04",x"96",x"F4",x"39",x"95",x"11",x"98",x"5F",x"C3",x"F2",x"C3",x"BE",x"0F",x"84",x"35",x"AF",x"15",x"91",x"F3",x"B3",x"39",x"EB",x"E6",x"D7",x"18",x"F0",x"90",x"DA",x"44",x"2E",x"65",x"6D",x"AC",x"6C",x"20",x"C8",x"60",x"F7",x"48",x"F3",x"CF",x"98",x"18",x"6D",x"F1",x"1F",x"A8",x"DB",x"C2",x"43",x"CA",x"70",x"49",x"99",x"38",x"94",x"56",x"8D",x"39",x"16",x"FB",x"5A",x"68",x"8A",x"29",x"CE",x"75",x"6F",x"09",x"C0",x"C2",x"40",x"18",x"60",x"6D",x"93",x"E0",x"EE",x"6E",x"C2",x"FE",x"EF",x"82",x"98",x"28",x"C2",x"2E",x"A5",x"D8",x"A5",x"13",x"60",x"EE",x"17",x"AD",x"59",x"F0",x"B2",x"F8",x"11",x"10",x"9A",x"D6",x"61",x"14",x"5C",x"0A",x"54",x"4A",x"5C",x"55",x"0E",x"99",x"6B",x"5E",x"CC",x"F9",x"18",x"F3",x"E0",x"61",x"96",x"6D",x"82",x"52",x"56",x"6E",x"0F",x"2E",x"66",x"DC",x"01",x"C0",x"02",x"E2",x"47",x"61",x"D6",x"D0",x"99",x"60",x"9A",x"F1",x"28",x"F0",x"02",x"48",x"EB",x"5B",x"FA",x"A8",x"8A",x"19",x"2C",x"5C",x"B4",x"4A",x"19",x"F0",x"B5",x"10",x"85",x"FC",x"20",x"FF",x"FC",x"18",x"B0",x"09",x"AE",x"37",x"FF",x"D9",x"65",x"55",x"E3",x"4E",x"FC",x"F7",x"66",x"51",x"94",x"CF",x"7D",x"08",x"20",x"13",x"5C",x"B0",x"05",x"4C",x"01",x"19",x"FA",x"BB",x"24",x"8C",x"9E",x"20",x"85",x"1F",x"10",x"C8",x"0B",x"D2",x"60",x"90",x"AD",x"E2",x"71",x"FB",x"A8",x"ED",x"69",x"19",x"4A",x"D5",x"34",x"E4",x"01",x"5E",x"20",x"A5",x"AD",x"68",x"A8",x"64",x"AF",x"94",x"FF",x"4D",x"65",x"95",x"2D",x"15",x"36",x"15",x"D7",x"C2",x"E8",x"62",x"17",x"84",x"0D",x"3C",x"4C",x"64",x"DC",x"19",x"AD",x"C3",x"DA",x"CD",x"BC",x"80",x"0A",x"20",x"AE",x"09",x"86",x"25",x"51",x"30",x"B2",x"32",x"92",x"89",x"D5",x"5A",x"37",x"C8",x"AB",x"66",x"80",x"36",x"EC",x"35",x"B1",x"54",x"EA",x"D9",x"2B",x"06",x"7A",x"71",x"93",x"18",x"E9",x"E8",x"8C",x"B0",x"1D",x"78",x"A9",x"41",x"3A",x"CB",x"63",x"00",x"26",x"B5",x"02",x"9F",x"D5",x"2A",x"20",x"E7",x"17",x"8C",x"FA",x"DF",x"33",x"3A",x"AA",x"61",x"7D",x"33",x"B1",x"FB",x"99",x"85",x"AC",x"B2",x"65",x"91",x"A5",x"9D",x"7B",x"FF",x"EE",x"34",x"3B",x"35",x"4B",x"BA",x"E8",x"AC",x"36",x"16",x"F3",x"18",x"76",x"C1",x"A7",x"05",x"45",x"D6",x"02",x"5A",x"46",x"87",x"31",x"C5",x"2D",x"48",x"CB",x"D0",x"1E",x"61",x"E4",x"C3",x"6A",x"0B",x"BD",x"C6",x"10",x"D3",x"14",x"F6",x"4C",x"1A",x"EC",x"22",x"36",x"1C",x"13",x"FD",x"1D",x"B2",x"58",x"92",x"F0",x"FD",x"68",x"F6",x"A5",x"42",x"B6",x"9E",x"C6",x"97",x"6C",x"11",x"ED",x"1A",x"58",x"B6",x"06",x"2C",x"1B",x"CB",x"56",x"71",x"81",x"1B",x"A6",x"B2",x"E0",x"9B",x"3F",x"4F",x"61",x"95",x"5C",x"7B",x"AB",x"0E",x"95",x"95",x"62",x"07",x"4D",x"D0",x"3D",x"A6",x"EF",x"1B",x"DA",x"37",x"0F",x"A2",x"CD",x"99",x"59",x"D0",x"20",x"20",x"CF",x"2C",x"2C",x"B9",x"B9",x"B7",x"17",x"15",x"B7",x"DE",x"F8",x"C3",x"B2",x"04",x"A3",x"3E",x"A0",x"C3",x"65",x"04",x"03",x"F2",x"F2",x"D3",x"44",x"4E",x"5C",x"80",x"26",x"1C",x"B8",x"D4",x"D3",x"53",x"06",x"E5",x"DD",x"EE",x"28",x"6A",x"51",x"67",x"65",x"43",x"60",x"16",x"83",x"37",x"80",x"78",x"F0",x"18",x"B9",x"35",x"60",x"1A",x"8D",x"8F",x"5D",x"A8",x"72",x"8F",x"45",x"20",x"C1",x"04",x"07",x"2B",x"06",x"10",x"BF",x"0B",x"10",x"4C",x"C0",x"4A",x"C6",x"A0",x"60",x"17",x"D0",x"D1",x"11",x"F8",x"56",x"05",x"E8",x"02",x"B5",x"6B",x"1D",x"BA",x"20",x"C1",x"2D",x"B0",x"F2",x"36",x"5B",x"EF",x"85",x"B4",x"A0",x"F9",x"08",x"E4",x"82",x"78",x"D5",x"F8",x"5D",x"34",x"81",x"DA",x"44",x"6C",x"13",x"39",x"55",x"02",x"16",x"1B",x"44",x"E4",x"C1",x"23",x"1F",x"9C",x"91",x"24",x"8E",x"1E",x"7C",x"0F",x"D9",x"E8",x"48",x"DC",x"32",x"71",x"20",x"36",x"3A",x"FD",x"D3",x"A2",x"AD",x"BE",x"09",x"EC",x"0A",x"1C",x"28",x"02",x"CB",x"50",x"62",x"CC",x"0F",x"08",x"D6",x"89",x"77",x"1D",x"70",x"5C",x"0C",x"A5",x"3D",x"05",x"69",x"9B",x"46",x"4C",x"26",x"1D",x"F3",x"31",x"4A",x"D9",x"B0",x"2D",x"5B",x"55",x"0A",x"B2",x"65",x"AD",x"B3",x"AA",x"C3",x"DD",x"30",x"1C",x"90",x"F6",x"02",x"80",x"18",x"4F",x"AE",x"14",x"10",x"9C",x"49",x"56",x"02",x"2D",x"06",x"48",x"A7",x"C9",x"34",x"B0",x"04",x"68",x"10",x"FF",x"1C",x"4B",x"5B",x"36",x"AA",x"02",x"7C",x"2F",x"6C",x"8A",x"A8",x"D4",x"28",x"A5",x"4C",x"21",x"1A",x"36",x"0D",x"16",x"52",x"BE",x"99",x"6D",x"F2",x"CA",x"86",x"29",x"DA",x"D0",x"20",x"ED",x"24",x"1C",x"19",x"DB",x"5D",x"C1",x"06",x"A4",x"B2",x"5D",x"73",x"81",x"D3",x"A8",x"95",x"1C",x"AD",x"DF",x"C0",x"02",x"EA",x"DB",x"AA",x"20",x"50",x"1D",x"80",x"D6",x"7F",x"14",x"BE",x"0D",x"77",x"0B",x"83",x"F0",x"C1",x"90",x"C0",x"46",x"12",x"9C",x"E4",x"05",x"4E",x"60",x"36",x"AF",x"09",x"68",x"54",x"10",x"1A",x"02",x"45",x"C9",x"20",x"34",x"14",x"16",x"69",x"47",x"A1",x"55",x"A1",x"17",x"51",x"0F",x"62",x"04",x"51",x"42",x"80",x"0D",x"70",x"03",x"3C",x"91",x"0D",x"98",x"29",x"48",x"80",x"9B",x"64",x"24",x"29",x"C7",x"3F",x"BA",x"F9",x"9C",x"74",x"CE",x"D3",x"E7",x"8E",x"D2",x"09",x"40",x"F8",x"10",x"A0",x"02",x"D6",x"5B",x"81",x"C0",x"21",x"1B",x"88",x"0C",x"A2",x"80",x"84",x"18",x"08",x"B2",x"56",x"29",x"BF",x"EA",x"E9",x"92",x"F7",x"20",x"9E",x"1D",x"A3",x"7F",x"0C",x"28",x"7E",x"00",x"56",x"7E",x"42",x"BD",x"72",x"D5",x"33",x"89",x"4A",x"75",x"37",x"CA",x"58",x"1E",x"AA",x"79",x"30",x"1A",x"AD",x"3A",x"75",x"0F",x"D7",x"E8",x"F8",x"12",x"C9",x"67",x"B0",x"0E",x"FC",x"37",x"6B",x"10",x"26",x"5F",x"CB",x"FC",x"1E",x"89",x"B7",x"1F",x"10",x"01",x"05",x"5A",x"18",x"FB",x"15",x"7A",x"7D",x"99",x"E7",x"A2",x"66",x"3E",x"4C",x"6B",x"1E",x"0F",x"E5",x"93",x"AD",x"30",x"46",x"02",x"B8",x"10",x"48",x"09",x"02",x"AA",x"71",x"5C",x"AA",x"4A",x"E9",x"D6",x"4F",x"32",x"59",x"0D",x"60",x"4F",x"2D",x"C6",x"B3",x"75",x"92",x"22",x"0E",x"9B",x"F7",x"C0",x"27",x"2D",x"7A",x"5C",x"02",x"71",x"1B",x"35",x"40",x"CD",x"68",x"16",x"93",x"F8",x"44",x"40",x"0F",x"80",x"0C",x"C6",x"65",x"8E",x"B3",x"58",x"6E",x"6A",x"02",x"60",x"E9",x"91",x"1E",x"41",x"56",x"9C",x"17",x"8C",x"31",x"8A",x"D3",x"4B",x"17",x"50",x"B3",x"F0",x"06",x"EE",x"1D",x"75",x"4C",x"1C",x"5A",x"30",x"F4",x"1F",x"ED",x"D8",x"38",x"F0",x"B6",x"09",x"3C",x"13",x"B3",x"A5",x"B2",x"E7",x"C9",x"06",x"F0",x"08",x"5F",x"02",x"0F",x"4C",x"45",x"1F",x"F9",x"58",x"52",x"AC",x"44",x"A8",x"C0",x"82",x"98",x"20",x"2D",x"20",x"46",x"AD",x"24",x"1B",x"25",x"8D",x"D1",x"2C",x"92",x"41",x"45",x"0D",x"BB",x"58",x"2F",x"0F",x"E6",x"B3",x"6E",x"B4",x"65",x"CA",x"D0",x"59",x"02",x"49",x"14",x"E3",x"2A",x"DE",x"43",x"E3",x"74",x"59",x"E2",x"80",x"B0",x"F3",x"B9",x"13",x"1F",x"3A",x"E4",x"95",x"AD",x"F0",x"B3",x"A2",x"C6",x"B8",x"79",x"CC",x"87",x"DE",x"F8",x"E6",x"AC",x"B6",x"68",x"A3",x"49",x"69",x"CA",x"D8",x"C2",x"68",x"52",x"1A",x"D2",x"B6",x"90",x"32",x"A6",x"3E",x"F0",x"ED",x"35",x"9F",x"BD",x"C1",x"DC",x"8F",x"C6",x"AC",x"58",x"B4",x"11",x"44",x"AA",x"A2",x"46",x"CF",x"A8",x"5B",x"4C",x"A3",x"C9",x"C4",x"7B",x"A5",x"2A",x"E9",x"A3",x"6A",x"8F",x"AA",x"A9",x"D1",x"A0",x"91",x"A8",x"B7",x"50",x"A7",x"52",x"B5",x"A5",x"0E",x"B6",x"30",x"10",x"D6",x"1E",x"BE",x"29",x"25",x"AE",x"39",x"0F",x"E2",x"1F",x"0F",x"49",x"58",x"18",x"69",x"01",x"74",x"80",x"0A",x"A6",x"A4",x"85",x"1A",x"15",x"99",x"52",x"DD",x"94",x"16",x"AD",x"53",x"27",x"FE",x"DB",x"72",x"0D",x"B0",x"55",x"34",x"3A",x"16",x"75",x"00",x"A6",x"F0",x"5B",x"B6",x"D9",x"18",x"A9",x"82",x"96",x"03",x"21",x"76",x"FF",x"55",x"A5",x"47",x"6D",x"4D",x"57",x"00",x"0F",x"41",x"BB",x"2A",x"65",x"7D",x"9D",x"35",x"51",x"42",x"3B",x"46",x"B4",x"01",x"44",x"FE",x"AB",x"D1",x"06",x"90",x"AE",x"0E",x"AE",x"0B",x"EC",x"12",x"D0",x"F0",x"FB",x"FB",x"3B",x"E1",x"B3",x"72",x"60",x"B4",x"A6",x"B7",x"1C",x"80",x"C1",x"20",x"AD",x"E7",x"C7",x"55",x"2A",x"70",x"07",x"B0",x"09",x"3E",x"40",x"D6",x"EA",x"36",x"67",x"20",x"B8",x"62",x"78",x"05",x"C8",x"C9",x"BC",x"CA",x"57",x"54",x"CB",x"57",x"89",x"0B",x"A8",x"9A",x"6A",x"42",x"8D",x"CF",x"D6",x"4C",x"F6",x"FD",x"6A",x"2F",x"B8",x"05",x"94",x"11",x"12",x"07",x"AD",x"1E",x"14",x"E8",x"3A",x"16",x"D4",x"A1",x"39",x"08",x"DA",x"1B",x"DA",x"92",x"BA",x"0C",x"B8",x"0A",x"14",x"07",x"18",x"20",x"F6",x"17",x"D0",x"FD",x"5B",x"28",x"FF",x"BA",x"85",x"46",x"1F",x"9F",x"46",x"0D",x"A2",x"A8",x"F3",x"21",x"E1",x"1D",x"C2",x"47",x"C3",x"28",x"71",x"C3",x"61",x"9B",x"F5",x"4F",x"36",x"00",x"96",x"B0",x"F3",x"20",x"01",x"27",x"DA",x"21",x"F9",x"02",x"4E",x"32",x"03",x"CD",x"2E",x"79",x"48",x"68",x"58",x"96",x"27",x"71",x"A7",x"7A",x"82",x"22",x"83",x"DE",x"18",x"54",x"0E",x"9C",x"45",x"0C",x"B8",x"0E",x"06",x"23",x"6D",x"70",x"0F",x"66",x"06",x"E0",x"0E",x"E1",x"1B",x"02",x"AA",x"04",x"0E",x"3C",x"14",x"4C",x"02",x"70",x"99",x"26",x"14",x"E0",x"1A",x"61",x"04",x"B4",x"10",x"CE",x"0C",x"1A",x"3C",x"21",x"8C",x"31",x"C0",x"A2",x"A2",x"01",x"4B",x"61",x"B8",x"A0",x"24",x"C1",x"2E",x"6A",x"06",x"C0",x"9E",x"28",x"D0",x"F9",x"6F",x"31",x"48",x"B5",x"01",x"49",x"D6",x"45",x"3A",x"72",x"A9",x"11",x"85",x"B1",x"77",x"7D",x"7D",x"48",x"B9",x"96",x"2A",x"6F",x"AD",x"C7",x"7A",x"CD",x"59",x"93",x"D0",x"ED",x"12",x"2D",x"0A",x"B0",x"A3",x"2A",x"0E",x"B1",x"55",x"40",x"07",x"CD",x"14",x"F0",x"96",x"E7",x"52",x"34",x"07",x"24",x"B2",x"3F",x"34",x"64",x"C5",x"98",x"79",x"3C",x"23",x"B3",x"38",x"15",x"CC",x"26",x"F9",x"A2",x"0D",x"38",x"BC",x"43",x"60",x"E0",x"8F",x"0A",x"60",x"A8",x"4F",x"57",x"29",x"49",x"AA",x"40",x"03",x"05",x"E4",x"00",x"AE",x"4B",x"EF",x"98",x"25",x"4C",x"32",x"17",x"A2",x"02",x"4A",x"72",x"D4",x"19",x"44",x"6A",x"36",x"65",x"92",x"A6",x"21",x"EF",x"DB",x"00",x"8D",x"25",x"D3",x"99",x"23",x"B7",x"AF",x"D7",x"D6",x"04",x"B0",x"7B",x"DD",x"0B",x"A5",x"96",x"29",x"58",x"C9",x"19",x"90",x"76",x"20",x"75",x"D4",x"24",x"83",x"E1",x"A1",x"F9",x"76",x"8D",x"24",x"9A",x"18",x"25",x"9A",x"92",x"92",x"6E",x"1D",x"CE",x"19",x"39",x"15",x"09",x"11",x"9A",x"A8",x"CA",x"B7",x"73",x"D0",x"F8",x"5C",x"98",x"AC",x"5A",x"CE",x"8A",x"48",x"6E",x"A6",x"7F",x"E0",x"D7",x"CE",x"DE",x"03",x"7A",x"36",x"7C",x"70",x"2B",x"28",x"B7",x"24",x"0D",x"F0",x"D0",x"25",x"E2",x"AD",x"AC",x"22",x"34",x"B7",x"3B",x"C9",x"21",x"A4",x"30",x"3D",x"4C",x"A9",x"23",x"77",x"10",x"DA",x"69",x"57",x"25",x"CF",x"08",x"08",x"00",x"67",x"0F",x"71",x"01",x"16",x"15",x"02",x"67",x"1B",x"71",x"03",x"12",x"22",x"B0",x"62",x"56",x"04",x"25",x"C9",x"24",x"90",x"17",x"A9",x"EA",x"05",x"4C",x"63",x"24",x"60",x"C5",x"FF",x"F0",x"1D",x"D0",x"BF",x"2A",x"61",x"29",x"AD",x"AE",x"22",x"78",x"25",x"BD",x"77",x"B4",x"75",x"C2",x"C9",x"A0",x"D7",x"CB",x"2F",x"C7",x"24",x"B5",x"5B",x"73",x"ED",x"20",x"8D",x"27",x"2E",x"89",x"4A",x"06",x"EB",x"33",x"20",x"C3",x"80",x"62",x"86",x"E9",x"20",x"32",x"21",x"74",x"8B",x"C7",x"41",x"49",x"90",x"EF",x"A2",x"54",x"45",x"E0",x"C4",x"05",x"23",x"19",x"29",x"E5",x"D2",x"03",x"4E",x"49",x"CA",x"86",x"48",x"5F",x"33",x"58",x"85",x"E8",x"2B",x"A0",x"D0",x"B7",x"00",x"37",x"01",x"E0",x"4E",x"21",x"10",x"E0",x"B2",x"53",x"7E",x"D3",x"DF",x"86",x"04",x"48",x"CA",x"DB",x"02",x"A2",x"13",x"7A",x"10",x"82",x"0C",x"33",x"2B",x"AE",x"2C",x"04",x"9A",x"49",x"E2",x"97",x"DB",x"7C",x"0D",x"C0",x"12",x"46",x"C6",x"8E",x"B1",x"0C",x"AC",x"50",x"A7",x"6E",x"E7",x"89",x"BB",x"33",x"B8",x"C7",x"30",x"19",x"AC",x"11",x"73",x"09",x"E5",x"D2",x"C5",x"8A",x"1D",x"F1",x"25",x"E4",x"5D",x"3B",x"20",x"D8",x"26",x"A4",x"F2",x"06",x"00",x"0F",x"1C",x"F6",x"F3",x"A0",x"C0",x"B1",x"AA",x"D7",x"B4",x"F5",x"C7",x"00",x"70",x"73",x"53",x"C0",x"3E",x"78",x"1F",x"70",x"8C",x"00",x"76",x"05",x"88",x"27",x"98",x"59",x"2A",x"4D",x"81",x"03",x"84",x"06",x"48",x"16",x"23",x"34",x"18",x"B2",x"B4",x"B3",x"75",x"C1",x"FC",x"51",x"14",x"8B",x"A5",x"A7",x"D0",x"1F",x"83",x"B3",x"F0",x"01",x"67",x"85",x"95",x"5D",x"91",x"A8",x"60",x"B8",x"3D",x"0A",x"A3",x"99",x"01",x"24",x"03",x"96",x"DE",x"38",x"8B",x"BC",x"85",x"AD",x"B1",x"44",x"B8",x"E6",x"87",x"A2",x"D4",x"5C",x"F0",x"06",x"C8",x"E8",x"E4",x"AD",x"D0",x"FE",x"F6",x"86",x"8C",x"57",x"1A",x"FB",x"E2",x"0E",x"AA",x"11",x"96",x"AB",x"35",x"46",x"27",x"BF",x"E5",x"AD",x"4F",x"65",x"AC",x"8D",x"77",x"A5",x"42",x"CB",x"04",x"95",x"6D",x"45",x"D0",x"A8",x"A9",x"6B",x"02",x"E8",x"44",x"A7",x"C3",x"D9",x"A5",x"B3",x"A3",x"CE",x"88",x"48",x"B4",x"0D",x"F3",x"07",x"20",x"90",x"47",x"BE",x"F3",x"B9",x"00",x"4A",x"C4",x"FC",x"94",x"5C",x"FE",x"8E",x"68",x"48",x"11",x"3D",x"B3",x"F4",x"A6",x"47",x"67",x"44",x"AA",x"18",x"76",x"9D",x"25",x"05",x"A5",x"96",x"B1",x"07",x"F6",x"0F",x"3F",x"51",x"77",x"A4",x"4C",x"90",x"84",x"27",x"8B",x"54",x"75",x"D1",x"48",x"DF",x"22",x"61",x"68",x"97",x"28",x"16",x"DD",x"60",x"FE",x"48",x"19",x"6C",x"A7",x"92",x"8B",x"30",x"D3",x"BD",x"21",x"A9",x"DA",x"29",x"B6",x"00",x"30",x"B5",x"32",x"9E",x"7A",x"A0",x"FF",x"84",x"42",x"7E",x"E7",x"0A",x"A8",x"36",x"40",x"48",x"4C",x"12",x"B0",x"99",x"5D",x"DD",x"02",x"FD",x"A9",x"CC",x"37",x"40",x"7B",x"78",x"7B",x"76",x"84",x"44",x"C7",x"7C",x"6E",x"77",x"24",x"49",x"EA",x"29",x"90",x"03",x"4C",x"5B",x"28",x"18",x"FE",x"98",x"65",x"87",x"35",x"E2",x"04",x"4A",x"44",x"DD",x"5A",x"D0",x"E7",x"4C",x"CA",x"27",x"5D",x"E5",x"E0",x"14",x"DF",x"9B",x"C3",x"55",x"E8",x"4C",x"F6",x"27",x"F1",x"45",x"B5",x"05",x"8E",x"16",x"52",x"79",x"02",x"B5",x"06",x"94",x"D6",x"41",x"7B",x"01",x"57",x"35",x"A2",x"2B",x"EA",x"09",x"0A",x"C2",x"1E",x"AD",x"54",x"3B",x"50",x"46",x"0F",x"02",x"2B",x"53",x"96",x"61",x"1E",x"01",x"85",x"47",x"EE",x"29",x"56",x"20",x"6C",x"6A",x"89",x"E1",x"4C",x"4F",x"28",x"3F",x"3B",x"3D",x"F6",x"EB",x"16",x"17",x"0B",x"86",x"42",x"DE",x"F4",x"9D",x"65",x"31",x"DC",x"4B",x"A8",x"25",x"C7",x"0A",x"8D",x"AE",x"F1",x"00",x"22",x"ED",x"0D",x"04",x"4C",x"74",x"28",x"ED",x"2D",x"75",x"F4",x"A9",x"0C",x"FA",x"41",x"4B",x"A9",x"03",x"9D",x"84",x"43",x"8A",x"A8",x"4F",x"F0",x"13",x"F6",x"6A",x"B1",x"40",x"D2",x"AA",x"CA",x"DD",x"A4",x"43",x"B9",x"C8",x"92",x"4C",x"78",x"28",x"7F",x"8D",x"5E",x"5B",x"43",x"3E",x"60",x"A6",x"46",x"71",x"DB",x"BA",x"28",x"A6",x"F0",x"32",x"78",x"18",x"02",x"54",x"63",x"A0",x"35",x"B5",x"21",x"69",x"D0",x"A8",x"AD",x"88",x"9A",x"04",x"B6",x"81",x"90",x"21",x"49",x"D3",x"D4",x"08",x"C3",x"4B",x"4C",x"30",x"29",x"E0",x"06",x"D0",x"1D",x"FE",x"EB",x"75",x"09",x"04",x"4E",x"48",x"2C",x"EA",x"FB",x"A9",x"0A",x"E8",x"1D",x"F1",x"48",x"20",x"2A",x"B3",x"06",x"AA",x"A2",x"FF",x"60",x"E8",x"49",x"F5",x"30",x"E7",x"CE",x"A5",x"BA",x"DA",x"76",x"EB",x"14",x"E5",x"07",x"60",x"5F",x"76",x"A9",x"14",x"43",x"FB",x"C5",x"5A",x"FC",x"C8",x"91",x"97",x"18",x"A9",x"02",x"65",x"3E",x"34",x"FD",x"A5",x"3D",x"FE",x"9A",x"0C",x"DE",x"A5",x"E1",x"83",x"8B",x"AE",x"39",x"89",x"68",x"BD",x"1E",x"30",x"A4",x"50",x"F5",x"29",x"A6",x"40",x"CE",x"D9",x"5E",x"E2",x"A9",x"FF",x"26",x"1A",x"50",x"EA",x"24",x"94",x"2A",x"97",x"4D",x"87",x"64",x"2B",x"51",x"DC",x"70",x"D0",x"04",x"3B",x"36",x"2E",x"51",x"EA",x"F8",x"9E",x"9F",x"E5",x"60",x"6A",x"C8",x"8A",x"48",x"9C",x"2A",x"16",x"01",x"43",x"29",x"28",x"48",x"49",x"01",x"FA",x"44",x"10",x"41",x"1A",x"84",x"05",x"B1",x"BF",x"2F",x"49",x"1C",x"2F",x"12",x"87",x"8A",x"6B",x"02",x"1E",x"13",x"11",x"68",x"10",x"95",x"AA",x"E8",x"8E",x"B9",x"02",x"D9",x"2D",x"ED",x"85",x"65",x"05",x"43",x"0E",x"A0",x"29",x"17",x"16",x"F0",x"1F",x"30",x"2A",x"09",x"28",x"4C",x"FE",x"A0",x"4E",x"10",x"B1",x"DD",x"1E",x"30",x"5B",x"34",x"6D",x"DC",x"69",x"A8",x"13",x"16",x"60",x"12",x"DD",x"01",x"16",x"6D",x"A4",x"1F",x"58",x"01",x"11",x"4C",x"12",x"C0",x"C7",x"7A",x"50",x"4C",x"06",x"50",x"9A",x"A9",x"2D",x"84",x"C5",x"A4",x"C0",x"AE",x"91",x"C6",x"1A",x"58",x"2B",x"D1",x"93",x"1C",x"E4",x"4D",x"22",x"8A",x"04",x"25",x"C9",x"30",x"8E",x"38",x"E9",x"09",x"FE",x"1F",x"80",x"09",x"75",x"07",x"1F",x"9D",x"90",x"15",x"A2",x"60",x"0B",x"A2",x"21",x"64",x"65",x"AF",x"48",x"66",x"74",x"8D",x"C5",x"67",x"C3",x"1E",x"20",x"9E",x"61",x"59",x"D3",x"81",x"E3",x"30",x"0B",x"E5",x"AC",x"60",x"D0",x"09",x"E4",x"B2",x"F8",x"F0",x"0A",x"64",x"57",x"30",x"05",x"BD",x"E9",x"5E",x"71",x"59",x"E8",x"70",x"72",x"FD",x"41",x"6F",x"8F",x"0B",x"C0",x"08",x"D8",x"DE",x"3A",x"6B",x"55",x"1E",x"55",x"38",x"00",x"9F",x"26",x"05",x"D0",x"AC",x"E7",x"6A",x"1E",x"E7",x"2D",x"46",x"00",x"91",x"39",x"0C",x"58",x"CF",x"39",x"64",x"2C",x"76",x"A5",x"20",x"ED",x"18",x"8E",x"13",x"24",x"59",x"60",x"60",x"8E",x"BE",x"E6",x"E0",x"3C",x"78",x"59",x"C6",x"52",x"8C",x"70",x"72",x"04",x"EE",x"75",x"67",x"08",x"64",x"FA",x"63",x"12",x"D1",x"66",x"65",x"62",x"02",x"9F",x"6A",x"25",x"01",x"1D",x"6C",x"07",x"6A",x"75",x"F6",x"4B",x"06",x"87",x"72",x"03",x"6D",x"61",x"79",x"05",x"FD",x"6E",x"45",x"76",x"11",x"6F",x"63",x"74",x"10",x"73",x"65",x"FF",x"70",x"5B",x"FF",x"04",x"03",x"07",x"AF",x"08",x"06",x"05",x"01",x"0B",x"FA",x"0A",x"09",x"02",x"72",x"67",x"E1",x"1A",x"1E",x"25",x"8C",x"40",x"1F",x"20",x"FF",x"3E",x"BD",x"08",x"23",x"30",x"90",x"31",x"69",x"C6",x"B7",x"71",x"FB",x"A9",x"99",x"1B",x"26",x"80",x"13",x"13",x"0F",x"44",x"74",x"90",x"0A",x"37",x"40",x"43",x"EC",x"40",x"EA",x"EE",x"35",x"B5",x"C9",x"02",x"2C",x"35",x"AE",x"CD",x"2E",x"05",x"A2",x"01",x"56",x"E7",x"10",x"8E",x"72",x"5A",x"CA",x"1B",x"29",x"03",x"F0",x"0D",x"0F",x"21",x"1D",x"52",x"28",x"C9",x"9D",x"91",x"72",x"C9",x"1E",x"90",x"F8",x"A9",x"29",x"BF",x"45",x"41",x"54",x"62",x"8C",x"5A",x"2D",x"65",x"54",x"6C",x"26",x"8D",x"6B",x"88",x"A3",x"31",x"AA",x"14",x"12",x"C9",x"0D",x"90",x"F7",x"B9",x"12",x"55",x"12",x"1D",x"7A",x"86",x"01",x"96",x"3F",x"39",x"B5",x"6C",x"ED",x"AC",x"A5",x"DA",x"8A",x"91",x"CD",x"A5",x"90",x"BC",x"0C",x"AE",x"1F",x"BB",x"35",x"C2",x"2C",x"71",x"5C",x"45",x"60",x"3A",x"02",x"FD",x"2D",x"8A",x"C9",x"40",x"0C",x"F7",x"F0",x"16",x"C9",x"A0",x"F7",x"B0",x"10",x"03",x"4A",x"A4",x"2A",x"6E",x"B9",x"CE",x"B5",x"C8",x"AA",x"80",x"02",x"A2",x"5A",x"AD",x"FC",x"66",x"C9",x"0A",x"B0",x"07",x"8A",x"18",x"6D",x"7F",x"AA",x"B2",x"60",x"95",x"09",x"5D",x"D6",x"43",x"F2",x"A2",x"1C",x"37",x"2D",x"9D",x"65",x"82",x"EB",x"FA",x"A6",x"B4",x"DD",x"1B",x"29",x"33",x"09",x"AB",x"B3",x"1E",x"F0",x"0E",x"FD",x"AA",x"B2",x"5F",x"81",x"A4",x"6E",x"3B",x"D0",x"F5",x"A4",x"B3",x"AD",x"7F",x"B2",x"99",x"F6",x"B4",x"04",x"22",x"EF",x"4F",x"70",x"1A",x"A6",x"64",x"DA",x"81",x"D9",x"B1",x"2C",x"F0",x"F2",x"02",x"80",x"0B",x"83",x"B7",x"83",x"5A",x"C8",x"C0",x"EA",x"7D",x"EB",x"FA",x"37",x"20",x"E8",x"88",x"C4",x"B3",x"D0",x"0E",x"7F",x"84",x"86",x"F1",x"CA",x"16",x"91",x"71",x"21",x"97",x"3F",x"BF",x"1B",x"C2",x"0C",x"D0",x"C6",x"38",x"FD",x"A1",x"1F",x"8F",x"CD",x"20",x"5E",x"2F",x"3B",x"3C",x"19",x"C8",x"A2",x"0C",x"DB",x"45",x"07",x"21",x"1E",x"8D",x"D7",x"CD",x"98",x"CA",x"D0",x"CB",x"FA",x"89",x"39",x"54",x"93",x"1C",x"41",x"D3",x"1E",x"88",x"D8",x"48",x"56",x"37",x"32",x"39",x"61",x"7A",x"78",x"60",x"95",x"78",x"04",x"5C",x"25",x"70",x"62",x"78",x"6E",x"A8",x"20",x"89",x"2D",x"5E",x"A4",x"5D",x"A0",x"9B",x"C8",x"5A",x"6F",x"23",x"A3",x"7A",x"F9",x"74",x"2C",x"F7",x"84",x"1B",x"E8",x"C2",x"E0",x"03",x"D0",x"EF",x"77",x"2D",x"CA",x"D3",x"61",x"47",x"AD",x"F4",x"8C",x"1C",x"8C",x"E0",x"CC",x"7A",x"AA",x"26",x"D0",x"05",x"AD",x"63",x"0D",x"91",x"FD",x"21",x"41",x"8D",x"6D",x"CF",x"20",x"35",x"2B",x"AC",x"7D",x"59",x"5A",x"25",x"86",x"5B",x"0A",x"4F",x"D4",x"C8",x"A6",x"DC",x"A5",x"AA",x"44",x"09",x"70",x"9D",x"B9",x"DF",x"E6",x"43",x"68",x"7B",x"69",x"03",x"A8",x"B7",x"AF",x"D8",x"98",x"10",x"5C",x"03",x"ED",x"1A",x"AB",x"A8",x"04",x"0A",x"8A",x"80",x"43",x"17",x"B6",x"0E",x"E4",x"14",x"AD",x"5C",x"08",x"DC",x"E7",x"E4",x"26",x"B9",x"E5",x"B6",x"4A",x"76",x"70",x"49",x"56",x"C9",x"1F",x"C1",x"5B",x"A0",x"4C",x"FC",x"DC",x"A9",x"D1",x"F5",x"6D",x"A0",x"98",x"A5",x"2A",x"9B",x"8E",x"8D",x"4D",x"C8",x"AA",x"CA",x"EC",x"E1",x"0C",x"8D",x"CB",x"52",x"AC",x"B6",x"AD",x"59",x"6C",x"09",x"E5",x"EE",x"58",x"2F",x"EE",x"C8",x"B2",x"A4",x"7E",x"E3",x"60",x"98",x"48",x"2F",x"9D",x"FA",x"D3",x"B9",x"B6",x"FC",x"D3",x"48",x"54",x"D4",x"BB",x"A6",x"44",x"06",x"D4",x"DE",x"68",x"01",x"B4",x"C9",x"7B",x"8D",x"28",x"FC",x"38",x"A9",x"28",x"E5",x"F9",x"4A",x"AF",x"18",x"65",x"8B",x"46",x"4A",x"A4",x"44",x"F0",x"4A",x"C7",x"EB",x"37",x"3A",x"4A",x"F4",x"34",x"B3",x"60",x"85",x"18",x"A0",x"0F",x"04",x"49",x"0A",x"C8",x"E9",x"EB",x"03",x"96",x"B0",x"F8",x"01",x"E2",x"87",x"AD",x"5A",x"6F",x"40",x"83",x"BB",x"AA",x"71",x"C0",x"4A",x"FA",x"29",x"02",x"53",x"04",x"F5",x"30",x"01",x"56",x"A9",x"7E",x"0C",x"F6",x"D7",x"AD",x"5E",x"AE",x"D0",x"0D",x"BA",x"87",x"42",x"08",x"4C",x"D1",x"AF",x"BE",x"DF",x"55",x"52",x"67",x"E0",x"30",x"A0",x"27",x"BE",x"5F",x"52",x"86",x"04",x"3A",x"87",x"7A",x"00",x"D7",x"2F",x"65",x"18",x"04",x"A5",x"28",x"88",x"D8",x"B9",x"FF",x"67",x"F4",x"31",x"0B",x"C1",x"08",x"B7",x"40",x"DE",x"DB",x"52",x"6B",x"CA",x"8B",x"34",x"01",x"90",x"E9",x"00",x"90",x"6B",x"AB",x"02",x"3A",x"20",x"8A",x"40",x"D0",x"03",x"3A",x"AD",x"B0",x"9B",x"21",x"41",x"9B",x"1B",x"F4",x"5B",x"D8",x"08",x"F4",x"70",x"04",x"35",x"64",x"40",x"61",x"D9",x"EF",x"DF",x"7B",x"B0",x"03",x"EB",x"38",x"E9",x"20",x"60",x"48",x"A6",x"42",x"7F",x"3D",x"0D",x"D6",x"C9",x"FF",x"F0",x"51",x"29",x"0F",x"6B",x"3F",x"01",x"4B",x"31",x"BD",x"02",x"D5",x"37",x"85",x"FC",x"BD",x"E7",x"FB",x"29",x"8C",x"10",x"AA",x"0F",x"B5",x"50",x"A6",x"88",x"6E",x"60",x"C7",x"FF",x"C9",x"70",x"F0",x"01",x"1E",x"C8",x"90",x"B1",x"FB",x"48",x"5F",x"42",x"FA",x"69",x"04",x"AA",x"7A",x"CF",x"15",x"4B",x"BD",x"E8",x"36",x"5D",x"64",x"18",x"C5",x"02",x"EA",x"04",x"62",x"8D",x"CB",x"FE",x"85",x"A6",x"16",x"A8",x"3A",x"68",x"91",x"A5",x"7A",x"C2",x"FB",x"82",x"ED",x"9F",x"B0",x"11",x"7A",x"47",x"09",x"53",x"C4",x"2F",x"6A",x"41",x"2C",x"58",x"10",x"7A",x"30",x"D0",x"82",x"D7",x"80",x"D6",x"D8",x"E9",x"7F",x"F5",x"2B",x"8E",x"63",x"DD",x"26",x"08",x"B3",x"5E",x"69",x"DC",x"24",x"2C",x"8D",x"0F",x"75",x"EA",x"CB",x"13",x"B6",x"42",x"03",x"DA",x"1A",x"18",x"D4",x"CA",x"8E",x"FD",x"2A",x"66",x"07",x"93",x"22",x"3F",x"EA",x"02",x"DD",x"BA",x"E5",x"01",x"D6",x"2F",x"85",x"D1",x"00",x"25",x"6B",x"04",x"40",x"BD",x"05",x"55",x"A9",x"81",x"BA",x"0D",x"9E",x"91",x"85",x"F9",x"11",x"D5",x"0E",x"A4",x"F0",x"3D",x"61",x"09",x"B8",x"7B",x"F8",x"60",x"DA",x"09",x"0B",x"3F",x"01",x"C7",x"F8",x"3E",x"83",x"D7",x"BA",x"83",x"B5",x"82",x"14",x"45",x"28",x"A3",x"08",x"C5",x"AA",x"52",x"C6",x"AF",x"9C",x"0C",x"2A",x"F1",x"4F",x"84",x"96",x"EF",x"40",x"31",x"38",x"21",x"A2",x"94",x"08",x"49",x"A1",x"2F",x"1F",x"10",x"C2",x"07",x"11",x"21",x"20",x"00",x"40",x"0A",x"CA",x"BB",x"55",x"D1",x"F4",x"AE",x"9B",x"DD",x"D7",x"DA",x"0B",x"AA",x"9E",x"33",x"13",x"F3",x"E4",x"EC",x"E0",x"5F",x"47",x"5F",x"39",x"4B",x"4F",x"D9",x"5B",x"02",x"15",x"62",x"CB",x"85",x"79",x"C7",x"81",x"FA",x"78",x"B5",x"D4",x"B8",x"CA",x"FE",x"8B",x"6F",x"F6",x"BD",x"63",x"32",x"9D",x"40",x"03",x"FD",x"E8",x"E0",x"B0",x"F5",x"AF",x"B9",x"27",x"94",x"90",x"0D",x"DA",x"F8",x"07",x"D4",x"AD",x"C5",x"26",x"15",x"D0",x"CC",x"A2",x"0F",x"0B",x"D7",x"A8",x"90",x"DC",x"A0",x"7B",x"B0",x"C0",x"EF",x"D0",x"E0",x"BD",x"A2",x"D1",x"5B",x"1B",x"6D",x"72",x"90",x"A0",x"EF",x"B0",x"C0",x"BD",x"D0",x"F7",x"E0",x"8A",x"60",x"D2",x"BD",x"2B",x"33",x"FB",x"80",x"7A",x"90",x"A0",x"EF",x"B0",x"C0",x"BD",x"63",x"AE",x"E0",x"2B",x"9D",x"54",x"D3",x"CA",x"10",x"AC",x"F5",x"29",x"B1",x"83",x"49",x"BC",x"4D",x"09",x"F0",x"EC",x"4B",x"2A",x"91",x"6B",x"D0",x"E5",x"ED",x"5A",x"FE",x"A5",x"33",x"CA",x"02",x"FF",x"7A",x"CE",x"2C",x"55",x"A9",x"86",x"7C",x"72",x"D0",x"1F",x"64",x"C2",x"11",x"AD",x"1B",x"D6",x"F6",x"F6",x"9E",x"83",x"99",x"76",x"60",x"D8",x"08",x"48",x"DA",x"5A",x"DB",x"A5",x"FF",x"47",x"D3",x"87",x"0F",x"2D",x"4E",x"32",x"4D",x"3C",x"CD",x"9A",x"D0",x"37",x"6C",x"5E",x"51",x"AB",x"80",x"8B",x"E1",x"78",x"0A",x"AA",x"72",x"81",x"15",x"53",x"BD",x"82",x"BD",x"85",x"AF",x"A0",x"1D",x"B1",x"FA",x"AE",x"20",x"0A",x"31",x"3F",x"73",x"99",x"C0",x"07",x"88",x"10",x"F3",x"EE",x"7F",x"61",x"2E",x"C9",x"B3",x"03",x"11",x"19",x"D3",x"87",x"09",x"38",x"9E",x"92",x"CA",x"68",x"60",x"F6",x"34",x"61",x"E9",x"B7",x"DB",x"61",x"0A",x"CE",x"25",x"D0",x"2D",x"DB",x"10",x"69",x"5E",x"DD",x"6E",x"56",x"08",x"AD",x"20",x"4B",x"15",x"07",x"51",x"0D",x"A5",x"A7",x"F0",x"17",x"AD",x"FC",x"C2",x"49",x"9A",x"3A",x"33",x"92",x"B1",x"65",x"29",x"7F",x"AE",x"5F",x"7D",x"51",x"09",x"80",x"91",x"A8",x"A0",x"00",x"7E",x"91",x"25",x"C3",x"AD",x"96",x"56",x"02",x"57",x"49",x"FF",x"8D",x"55",x"6F",x"06",x"CE",x"DA",x"03",x"45",x"8C",x"01",x"DC",x"26",x"AF",x"2F",x"19",x"ED",x"B9",x"82",x"E9",x"3C",x"78",x"47",x"CF",x"11",x"18",x"4A",x"76",x"A8",x"8A",x"6D",x"42",x"7B",x"79",x"ED",x"B9",x"65",x"4D",x"F3",x"4E",x"12",x"E1",x"BA",x"34",x"09",x"DD",x"ED",x"2D",x"51",x"9B",x"52",x"F7",x"41",x"42",x"DE",x"55",x"42",x"79",x"07",x"AD",x"1A",x"D4",x"47",x"62",x"6A",x"E9",x"02",x"29",x"7E",x"AC",x"7E",x"20",x"FE",x"35",x"EC",x"8C",x"3D",x"B3",x"90",x"52",x"0A",x"48",x"8A",x"2A",x"AA",x"FE",x"68",x"8D",x"1B",x"C1",x"31",x"45",x"A8",x"8E",x"9E",x"68",x"1C",x"F7",x"AA",x"CC",x"EE",x"ED",x"5B",x"10",x"09",x"76",x"4F",x"3D",x"50",x"D9",x"48",x"48",x"35",x"8A",x"CC",x"F7",x"ED",x"B7",x"30",x"06",x"AC",x"EC",x"53",x"AE",x"A7",x"54",x"8C",x"2B",x"A2",x"8E",x"B6",x"D1",x"8D",x"69",x"35",x"98",x"20",x"85",x"36",x"7E",x"16",x"8A",x"35",x"55",x"12",x"5D",x"5D",x"13",x"0D",x"DC",x"DE",x"FB",x"7A",x"FA",x"68",x"28",x"40",x"FF",x"24",x"45",x"B5",x"2C",x"CD",x"33",x"B6",x"B2",x"BC",x"CA",x"72",x"ED",x"74",x"95",x"05",x"47",x"45",x"4E",x"14",x"46",x"62",x"19",x"01",x"6B",x"42",x"F3",x"4A",x"41",x"DE",x"49",x"7B",x"B3",x"CB",x"3F",x"8C",x"56",x"29",x"9B",x"D0",x"08",x"ED",x"CD",x"19",x"F0",x"3A",x"DB",x"91",x"34",x"EE",x"ED",x"28",x"1A",x"0B",x"87",x"47",x"38",x"51",x"48",x"88",x"68",x"29",x"D3",x"80",x"59",x"4D",x"97",x"D0",x"B5",x"0F",x"44",x"EB",x"18",x"B0",x"43",x"AB",x"66",x"B2",x"4C",x"FD",x"35",x"EE",x"3E",x"F5",x"40",x"D2",x"8C",x"B4",x"C6",x"8D",x"42",x"ED",x"59",x"C6",x"82",x"3F",x"B0",x"EE",x"00",x"23",x"68",x"C9",x"C0",x"90",x"07",x"6F",x"A2",x"FF",x"C8",x"38",x"AC",x"A7",x"5A",x"8A",x"A7",x"18",x"60",x"0F",x"CD",x"49",x"33",x"20",x"A6",x"64",x"10",x"85",x"13",x"57",x"A3",x"21",x"D0",x"0C",x"B7",x"48",x"29",x"76",x"F0",x"05",x"A9",x"74",x"3D",x"58",x"7B",x"55",x"5B",x"56",x"56",x"49",x"9A",x"18",x"B7",x"4A",x"B8",x"64",x"30",x"AD",x"50",x"74",x"C9",x"00",x"F0",x"FB",x"88",x"09",x"01",x"C8",x"84",x"58",x"89",x"29",x"FE",x"5D",x"10",x"5B",x"18",x"B6",x"4B",x"96",x"8D",x"C6",x"2A",x"4C",x"56",x"69",x"94",x"35",x"5C",x"2A",x"AD",x"5B",x"32",x"8D",x"01",x"FA",x"D0",x"60",x"37",x"15",x"A0",x"04",x"F0",x"05",x"58",x"06",x"08",x"10",x"07",x"00",x"28",x"50",x"78",x"A0",x"C8",x"F0",x"FF",x"18",x"40",x"68",x"90",x"B8",x"E0",x"08",x"30",x"FF",x"58",x"80",x"A8",x"D0",x"F8",x"20",x"48",x"70",x"FF",x"98",x"C0",x"17",x"D8",x"1E",x"D9",x"0B",x"DA",x"01",x"DB",x"22",x"91",x"D0",x"78",x"38",x"B3",x"22",x"9A",x"99",x"88",x"D0",x"5E",x"85",x"BB",x"B3",x"22",x"22",x"1A",x"19",x"10",x"08",x"02",x"21",x"91",x"91",x"08",x"B9",x"84",x"22",x"99",x"E6",x"07",x"88",x"D0",x"F7",x"18",x"AA",x"98",x"29",x"0F",x"99",x"68",x"03",x"F0",x"0C",x"8A",x"79",x"67",x"03",x"99",x"68",x"03",x"A5",x"9F",x"79",x"9B",x"03",x"99",x"9C",x"03",x"A9",x"01",x"85",x"9F",x"A9",x"78",x"20",x"00",x"01",x"4A",x"AA",x"F0",x"09",x"08",x"06",x"9F",x"38",x"6A",x"CA",x"D0",x"F9",x"28",x"6A",x"99",x"34",x"03",x"30",x"05",x"A5",x"9F",x"86",x"9F",x"24",x"8A",x"C8",x"C0",x"34",x"D0",x"C1",x"A0",x"00",x"8A",x"4C",x"9C",x"01",x"22",x"00",x"37",x"69",x"80",x"0A",x"10",x"0F",x"06",x"FD",x"D0",x"08",x"48",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"68",x"2A",x"30",x"F1",x"70",x"01",x"60",x"38",x"85",x"A7",x"AD",x"29",x"01",x"D0",x"06",x"CE",x"2A",x"01",x"8E",x"E7",x"DB",x"CE",x"29",x"01",x"AD",x"8E",x"21",x"60",x"20",x"1A",x"01",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"66",x"A8",x"CA",x"06",x"FD",x"D0",x"06",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"E8",x"90",x"F3",x"F0",x"E1",x"E0",x"11",x"B0",x"51",x"BD",x"33",x"03",x"20",x"00",x"01",x"7D",x"67",x"03",x"85",x"9E",x"AA",x"24",x"A8",x"10",x"09",x"70",x"07",x"A9",x"00",x"20",x"05",x"01",x"D0",x"25",x"A9",x"F1",x"E0",x"03",x"B0",x"03",x"BD",x"A2",x"01",x"B8",x"20",x"05",x"01",x"18",x"AA",x"BD",x"34",x"03",x"20",x"00",x"01",x"7D",x"68",x"03",x"85",x"AE",x"A5",x"A7",x"7D",x"9C",x"03",x"65",x"FF",x"85",x"AF",x"A6",x"9E",x"B1",x"AE",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"CA",x"D0",x"F1",x"86",x"A7",x"F0",x"99",x"4C",x"0D",x"08",x"CC",x"F2",x"01",x"00",x"0B",x"08",x"0A",x"7C",x"9E",x"32",x"30",x"FA",x"31",x"53",x"A7",x"4C",x"47",x"11",x"5C",x"52",x"E8",x"50",x"53",x"09",x"C5",x"9A",x"2E",x"53",x"41",x"A4",x"A2",x"3D",x"43",x"4F",x"4E",x"46",x"49",x"FD",x"55",x"A8",x"52",x"45",x"20",x"4D",x"45",x"47",x"41",x"BF",x"71",x"B5",x"91",x"0C",x"6C",x"6A",x"27",x"50",x"52",x"4F",x"50",x"2E",x"4D",x"36",x"35",x"55",x"2E",x"4E",x"41",x"4D",x"45",x"3D",x"43",x"4F",x"4E",x"46",x"49",x"47",x"55",x"52",x"45",x"20",x"4D",x"45",x"47",x"41",x"36",x"35",x"4D",x"36",x"35",x"55",x"53",x"44",x"43",x"41",x"52",x"44",x"20",x"46",x"44",x"49",x"53",x"4B",x"2B",x"46",x"4F",x"52",x"4D",x"41",x"54",x"20",x"55",x"54",x"49",x"4C",x"49",x"54",x"59",x"00",x"00",x"00",x"00",x"00",x"91",x"33",x"0D",x"08",x"56",x"23",x"13",x"57",x"01",x"08",x"0B",x"08",x"37",x"01",x"9E",x"32",x"30",x"36",x"31",x"00",x"00",x"00",x"BA",x"BD",x"88",x"3A",x"9D",x"FC",x"00",x"CA",x"D0",x"F7",x"A0",x"35",x"4C",x"3A",x"3A",x"85",x"FF",x"90",x"94",x"EB",x"9A",x"AE",x"93",x"79",x"F4",x"86",x"01",x"60",x"63",x"57",x"16",x"0B",x"45",x"6C",x"B0",x"AA",x"C1",x"82",x"3B",x"33",x"00",x"3B",x"93",x"A2",x"BE",x"41",x"2E",x"50",x"D7",x"81",x"5E",x"18",x"E6",x"A0",x"05",x"E0",x"B1",x"93",x"83",x"F2",x"73",x"A9",x"19",x"4F",x"F0",x"0F",x"25",x"44",x"23",x"63",x"07",x"61",x"68",x"1A",x"AE",x"1C",x"D8",x"EE",x"7E",x"A8",x"22",x"33",x"7C",x"18",x"0D",x"AC",x"1F",x"43",x"ED",x"56",x"03",x"6A",x"03",x"36",x"FF",x"2D",x"24",x"61",x"3C",x"99",x"3E",x"33",x"68",x"18",x"79",x"58",x"17",x"EF",x"A8",x"F0",x"D7",x"E7",x"A0",x"E1",x"F4",x"C0",x"F3",x"F3",x"F2",x"F1",x"BC",x"37",x"F5",x"88",x"AE",x"F6",x"D2",x"7C",x"E2",x"D3",x"63",x"21",x"F8",x"0A",x"EB",x"F6",x"78",x"C0",x"3D",x"65",x"15",x"58",x"E3",x"E0",x"06",x"81",x"96",x"18",x"72",x"00",x"63",x"EF",x"83",x"3D",x"39",x"16",x"B8",x"77",x"08",x"18",x"99",x"81",x"07",x"0A",x"33",x"34",x"23",x"FA",x"57",x"69",x"61",x"02",x"12",x"F6",x"18",x"51",x"19",x"AC",x"8D",x"3D",x"E6",x"47",x"BA",x"02",x"D1",x"20",x"F4",x"82",x"28",x"A4",x"EE",x"47",x"76",x"86",x"F2",x"34",x"93",x"7B",x"75",x"89",x"76",x"71",x"D2",x"B9",x"16",x"E5",x"B4",x"25",x"00",x"18",x"E1",x"5C",x"02",x"18",x"64",x"B3",x"38",x"52",x"B9",x"A2",x"C3",x"C5",x"96",x"17",x"E4",x"5D",x"02",x"CA",x"28",x"F0",x"97",x"44",x"A0",x"2F",x"90",x"16",x"D0",x"92",x"20",x"21",x"40",x"05",x"3A",x"40",x"72",x"90",x"B4",x"80",x"06",x"4A",x"90",x"A1",x"0E",x"35",x"0F",x"30",x"54",x"03",x"96",x"EE",x"C1",x"50",x"87",x"9A",x"07",x"18",x"EA",x"01",x"70",x"F7",x"60",x"28",x"0B",x"C0",x"54",x"44",x"4D",x"04",x"31",x"60",x"5C",x"01",x"52",x"CC",x"D5",x"93",x"81",x"04",x"FA",x"4A",x"43",x"2F",x"4F",x"67",x"C7",x"A6",x"73",x"35",x"62",x"D6",x"21",x"79",x"41",x"DE",x"1E",x"20",x"AF",x"23",x"FA",x"76",x"92",x"C6",x"97",x"96",x"6B",x"1B",x"D4",x"0E",x"BA",x"BF",x"0F",x"98",x"1C",x"77",x"31",x"27",x"60",x"5C",x"CA",x"0E",x"3E",x"30",x"70",x"CB",x"0B",x"48",x"93",x"36",x"8D",x"00",x"F9",x"12",x"35",x"3E",x"53",x"E2",x"E7",x"C7",x"9D",x"4B",x"09",x"89",x"58",x"13",x"9A",x"BC",x"1D",x"03",x"49",x"0E",x"3C",x"DA",x"06",x"4F",x"12",x"72",x"76",x"27",x"7B",x"2F",x"F0",x"1B",x"DF",x"60",x"77",x"D1",x"17",x"B8",x"F4",x"C5",x"50",x"05",x"84",x"0A",x"92",x"47",x"5C",x"19",x"1C",x"0D",x"B6",x"49",x"B1",x"D0",x"14",x"5C",x"9C",x"6F",x"EB",x"06",x"4C",x"70",x"C1",x"0F",x"97",x"D5",x"35",x"4D",x"E4",x"0C",x"03",x"BA",x"2A",x"CC",x"0D",x"79",x"88",x"51",x"F2",x"3D",x"38",x"44",x"22",x"3C",x"39",x"A8",x"A6",x"D7",x"88",x"AA",x"10",x"FC",x"6A",x"25",x"0A",x"48",x"68",x"F0",x"FF",x"17",x"2E",x"DD",x"BB",x"06",x"7A",x"81",x"DA",x"E3",x"A2",x"F4",x"14",x"35",x"5F",x"8C",x"50",x"DF",x"A8",x"74",x"C4",x"A0",x"71",x"54",x"08",x"B2",x"AE",x"C8",x"AC",x"B6",x"73",x"F0",x"0D",x"29",x"F2",x"07",x"33",x"A5",x"21",x"31",x"7D",x"62",x"8D",x"E3",x"80",x"0C",x"ED",x"2A",x"AA",x"52",x"62",x"28",x"81",x"9F",x"F1",x"76",x"59",x"C9",x"9F",x"74",x"47",x"58",x"72",x"5D",x"14",x"78",x"94",x"30",x"8D",x"8F",x"7F",x"80",x"0F",x"AD",x"87",x"A6",x"06",x"6C",x"CC",x"69",x"6F",x"04",x"25",x"27",x"87",x"1B",x"37",x"25",x"8A",x"7E",x"77",x"CF",x"D0",x"02",x"80",x"FE",x"5F",x"26",x"91",x"DD",x"03",x"85",x"FF",x"FB",x"04",x"78",x"8C",x"B9",x"64",x"B3",x"B5",x"9E",x"4A",x"8B",x"C5",x"19",x"70",x"97",x"03",x"15",x"6A",x"56",x"EA",x"60",x"A7",x"E0",x"23",x"C9",x"01",x"AD",x"3F",x"2B",x"0D",x"3E",x"F1",x"CC",x"82",x"11",x"16",x"13",x"D7",x"85",x"74",x"9C",x"6D",x"08",x"26",x"1D",x"AA",x"AC",x"6C",x"CF",x"7F",x"1A",x"76",x"C5",x"FE",x"52",x"DF",x"E0",x"EF",x"E1",x"79",x"E2",x"DA",x"DE",x"D9",x"F3",x"D8",x"D7",x"BC",x"5D",x"21",x"08",x"0B",x"BE",x"1F",x"CA",x"78",x"70",x"E7",x"E8",x"DE",x"E9",x"B3",x"67",x"84",x"F1",x"21",x"81",x"BA",x"3D",x"E5",x"C1",x"D4",x"8D",x"48",x"2A",x"8E",x"6B",x"9A",x"8C",x"30",x"93",x"11",x"61",x"30",x"23",x"C0",x"D6",x"FF",x"67",x"71",x"9C",x"9D",x"BD",x"9E",x"67",x"CB",x"08",x"03",x"DB",x"06",x"4C",x"80",x"B2",x"12",x"83",x"CD",x"03",x"E2",x"94",x"3E",x"0C",x"13",x"4A",x"13",x"3B",x"50",x"E9",x"03",x"72",x"60",x"8D",x"37",x"EF",x"81",x"3E",x"8A",x"F4",x"0F",x"93",x"F6",x"EA",x"0B",x"9C",x"54",x"43",x"0B",x"67",x"C4",x"9C",x"0E",x"A5",x"CC",x"17",x"A8",x"F5",x"A9",x"AA",x"9E",x"F0",x"33",x"AB",x"07",x"9D",x"8D",x"F9",x"7B",x"C3",x"BE",x"09",x"59",x"A8",x"6B",x"C9",x"0D",x"F5",x"21",x"DE",x"53",x"30",x"2D",x"07",x"0F",x"96",x"D6",x"1B",x"8D",x"F7",x"F8",x"F8",x"F9",x"9E",x"38",x"9B",x"62",x"4F",x"E9",x"A5",x"FA",x"F9",x"9E",x"F8",x"E7",x"F7",x"AD",x"19",x"FE",x"E2",x"FD",x"79",x"FC",x"FB",x"DE",x"C3",x"79",x"68",x"88",x"3D",x"2E",x"B9",x"11",x"57",x"BF",x"11",x"CD",x"6D",x"AC",x"91",x"18",x"40",x"E3",x"20",x"71",x"42",x"E2",x"07",x"4C",x"5E",x"BD",x"DF",x"D8",x"6E",x"D6",x"01",x"F3",x"4E",x"81",x"5E",x"B6",x"18",x"44",x"E7",x"2F",x"A2",x"E0",x"08",x"F9",x"CF",x"11",x"E3",x"E4",x"EF",x"E5",x"D9",x"33",x"C2",x"2B",x"DA",x"07",x"4A",x"C0",x"0D",x"3A",x"DB",x"99",x"DC",x"F7",x"DD",x"A5",x"AC",x"DE",x"7C",x"73",x"A3",x"3D",x"A2",x"4F",x"A1",x"4C",x"91",x"A0",x"95",x"AC",x"EA",x"AD",x"3D",x"AE",x"7B",x"46",x"13",x"58",x"FB",x"A0",x"02",x"B0",x"B1",x"DE",x"B2",x"B3",x"67",x"84",x"06",x"B5",x"0F",x"AB",x"CC",x"1F",x"4F",x"A8",x"42",x"A5",x"DD",x"A6",x"53",x"C6",x"A7",x"94",x"BC",x"C0",x"0F",x"D5",x"D2",x"1B",x"8D",x"B4",x"B5",x"BE",x"B6",x"0C",x"E7",x"F9",x"B7",x"78",x"60",x"3C",x"6C",x"B5",x"82",x"07",x"8C",x"F3",x"11",x"1C",x"FA",x"8D",x"75",x"E0",x"DE",x"AA",x"1C",x"61",x"22",x"D2",x"A4",x"9E",x"17",x"F9",x"33",x"83",x"67",x"EB",x"7D",x"68",x"AD",x"CB",x"B7",x"69",x"12",x"A6",x"B6",x"6A",x"FE",x"CF",x"81",x"3C",x"14",x"8D",x"85",x"1F",x"8E",x"8A",x"86",x"23",x"8C",x"87",x"7B",x"0F",x"57",x"14",x"88",x"0F",x"8D",x"89",x"C5",x"87",x"8E",x"8A",x"E2",x"08",x"E3",x"8B",x"0B",x"5E",x"18",x"8C",x"45",x"42",x"0C",x"5B",x"71",x"0F",x"8D",x"75",x"C5",x"87",x"8E",x"76",x"E2",x"08",x"A3",x"CA",x"77",x"BE",x"82",x"36",x"23",x"78",x"66",x"61",x"8D",x"79",x"2E",x"8E",x"7A",x"CC",x"04",x"89",x"2D",x"A8",x"6D",x"95",x"44",x"7C",x"A5",x"1A",x"10",x"EE",x"CC",x"C0",x"1D",x"71",x"7F",x"77",x"D6",x"AF",x"85",x"E3",x"B5",x"C0",x"77",x"01",x"EA",x"53",x"01",x"20",x"3E",x"0B",x"68",x"49",x"01",x"96",x"66",x"E9",x"48",x"99",x"94",x"91",x"35",x"4F",x"43",x"24",x"18",x"D6",x"D5",x"01",x"8E",x"59",x"04",x"F2",x"8E",x"2C",x"02",x"7D",x"46",x"5A",x"CA",x"85",x"F1",x"DA",x"E2",x"7D",x"41",x"16",x"52",x"D9",x"61",x"E1",x"48",x"8F",x"72",x"A6",x"93",x"55",x"94",x"AA",x"41",x"B7",x"95",x"12",x"61",x"8D",x"96",x"7B",x"C8",x"7B",x"D8",x"39",x"A2",x"01",x"A9",x"F8",x"62",x"B7",x"C9",x"6D",x"A8",x"C6",x"1B",x"98",x"F1",x"91",x"2F",x"0C",x"7E",x"22",x"EB",x"06",x"60",x"0A",x"C2",x"A9",x"66",x"D1",x"CB",x"9B",x"09",x"58",x"C1",x"B1",x"03",x"9B",x"D6",x"55",x"5B",x"AD",x"A9",x"A9",x"AA",x"8D",x"AE",x"7B",x"4D",x"2F",x"3E",x"11",x"0C",x"90",x"93",x"2F",x"23",x"86",x"B1",x"01",x"81",x"15",x"E6",x"BF",x"8F",x"50",x"72",x"1E",x"9F",x"EE",x"AF",x"04",x"E5",x"0B",x"C1",x"47",x"2E",x"8E",x"3D",x"AE",x"06",x"12",x"18",x"72",x"8B",x"0C",x"9E",x"E8",x"61",x"10",x"F6",x"57",x"87",x"7B",x"80",x"C0",x"F0",x"71",x"FA",x"78",x"0F",x"EE",x"64",x"3B",x"35",x"7A",x"18",x"54",x"EC",x"60",x"0F",x"3C",x"0D",x"E8",x"E1",x"8D",x"60",x"C4",x"62",x"C1",x"41",x"11",x"6F",x"B9",x"01",x"56",x"40",x"1A",x"00",x"AF",x"0A",x"8F",x"43",x"84",x"60",x"A4",x"AF",x"90",x"53",x"82",x"8A",x"A0",x"C9",x"21",x"4A",x"04",x"A0",x"D5",x"81",x"C8",x"0F",x"8D",x"EB",x"0F",x"B4",x"F8",x"0B",x"8F",x"64",x"79",x"0A",x"FB",x"96",x"15",x"82",x"A2",x"08",x"5C",x"38",x"0D",x"66",x"07",x"94",x"9A",x"F4",x"8D",x"D2",x"1D",x"DE",x"61",x"07",x"2A",x"9C",x"68",x"62",x"25",x"AF",x"56",x"56",x"10",x"C9",x"A5",x"FF",x"7B",x"2B",x"9E",x"10",x"A0",x"A5",x"F0",x"B9",x"18",x"10",x"1A",x"67",x"C1",x"3B",x"21",x"6C",x"28",x"AD",x"2A",x"89",x"58",x"EF",x"AA",x"C9",x"F0",x"B2",x"C7",x"70",x"F6",x"2A",x"AD",x"E5",x"F5",x"AB",x"E9",x"AD",x"4A",x"EB",x"D4",x"EC",x"7B",x"ED",x"F6",x"8C",x"30",x"EE",x"D2",x"ED",x"F3",x"EC",x"EC",x"7A",x"EB",x"7C",x"1F",x"11",x"CC",x"0D",x"C6",x"8C",x"19",x"FC",x"31",x"F1",x"79",x"F2",x"F3",x"58",x"CF",x"F4",x"F4",x"7C",x"5C",x"86",x"71",x"CF",x"6B",x"25",x"30",x"C4",x"07",x"05",x"CB",x"4E",x"35",x"E1",x"78",x"E2",x"B9",x"B7",x"77",x"C3",x"59",x"00",x"7E",x"19",x"7F",x"53",x"64",x"32",x"93",x"70",x"18",x"16",x"85",x"FA",x"91",x"82",x"7B",x"78",x"87",x"C4",x"83",x"65",x"22",x"0E",x"23",x"AA",x"77",x"BF",x"10",x"AC",x"15",x"D2",x"69",x"0D",x"7E",x"14",x"67",x"04",x"18",x"F0",x"1C",x"E1",x"1E",x"C3",x"B0",x"14",x"A9",x"08",x"45",x"00",x"24",x"5B",x"9C",x"0E",x"F7",x"30",x"E3",x"16",x"08",x"78",x"40",x"C4",x"53",x"28",x"0F",x"9E",x"E7",x"E7",x"2C",x"A5",x"29",x"98",x"99",x"18",x"A9",x"2E",x"6D",x"4B",x"87",x"B5",x"12",x"23",x"AE",x"8B",x"17",x"13",x"EB",x"08",x"62",x"86",x"B0",x"11",x"F1",x"D0",x"18",x"7C",x"93",x"47",x"AD",x"64",x"A0",x"57",x"33",x"74",x"6E",x"14",x"E6",x"20",x"AF",x"A3",x"B0",x"EC",x"80",x"B1",x"AD",x"14",x"B2",x"A6",x"9C",x"B3",x"34",x"E5",x"43",x"B4",x"52",x"A9",x"41",x"B5",x"D7",x"B6",x"7B",x"B7",x"B8",x"EF",x"B9",x"95",x"8D",x"BA",x"79",x"7E",x"BE",x"D2",x"A2",x"73",x"6B",x"39",x"39",x"C1",x"BF",x"29",x"79",x"E9",x"00",x"59",x"0A",x"18",x"EB",x"01",x"8D",x"CF",x"79",x"60",x"FC",x"1F",x"71",x"FF",x"D6",x"3E",x"4F",x"B9",x"19",x"74",x"9A",x"2F",x"5E",x"51",x"E9",x"11",x"DC",x"BE",x"B8",x"8A",x"C4",x"AF",x"F1",x"41",x"1B",x"22",x"07",x"28",x"51",x"78",x"41",x"2D",x"07",x"03",x"4D",x"0E",x"1C",x"AC",x"B0",x"82",x"02",x"70",x"03",x"04",x"3E",x"03",x"1E",x"6C",x"01",x"06",x"F5",x"04",x"B1",x"07",x"81",x"05",x"8F",x"24",x"06",x"08",x"A7",x"49",x"02",x"EF",x"D6",x"7A",x"A7",x"CA",x"8A",x"06",x"9A",x"42",x"F0",x"04",x"D3",x"DE",x"52",x"29",x"C1",x"C5",x"69",x"8B",x"0B",x"2F",x"FC",x"B0",x"E9",x"50",x"A6",x"B5",x"C1",x"8C",x"8D",x"EC",x"94",x"F0",x"06",x"48",x"49",x"68",x"7B",x"7E",x"4C",x"95",x"A4",x"03",x"7C",x"E2",x"35",x"B1",x"80",x"91",x"6E",x"17",x"43",x"9B",x"CD",x"F0",x"05",x"B4",x"EE",x"0C",x"31",x"51",x"3C",x"06",x"B7",x"30",x"1A",x"61",x"C4",x"1C",x"12",x"DC",x"8A",x"3F",x"18",x"36",x"2C",x"86",x"C9",x"93",x"CB",x"29",x"80",x"CA",x"DD",x"56",x"A8",x"16",x"0A",x"5A",x"24",x"C2",x"14",x"87",x"17",x"28",x"F0",x"13",x"E1",x"05",x"2B",x"7C",x"12",x"D8",x"01",x"35",x"1F",x"0D",x"FA",x"65",x"48",x"42",x"F8",x"0F",x"B0",x"C5",x"F0",x"7A",x"46",x"D8",x"E2",x"0E",x"30",x"70",x"36",x"7A",x"BC",x"B8",x"49",x"8D",x"30",x"13",x"C1",x"30",x"0D",x"E1",x"C6",x"BC",x"05",x"8A",x"9A",x"04",x"47",x"25",x"ED",x"95",x"73",x"59",x"53",x"34",x"91",x"04",x"22",x"4A",x"E6",x"E7",x"BC",x"4F",x"50",x"A1",x"C5",x"C9",x"F2",x"A2",x"14",x"B2",x"4F",x"7E",x"A0",x"8E",x"66",x"7E",x"D7",x"99",x"62",x"B3",x"D0",x"56",x"0C",x"75",x"A2",x"B9",x"07",x"A8",x"32",x"55",x"6C",x"8F",x"AD",x"6D",x"BA",x"C9",x"B6",x"B6",x"4A",x"3E",x"71",x"AD",x"16",x"87",x"8A",x"E7",x"A1",x"D4",x"6B",x"C8",x"DA",x"04",x"B0",x"0C",x"B2",x"FC",x"E1",x"0E",x"1B",x"36",x"9B",x"EE",x"DF",x"E2",x"7A",x"A2",x"62",x"AE",x"29",x"D6",x"8D",x"2E",x"AD",x"79",x"77",x"EC",x"81",x"EE",x"06",x"C9",x"82",x"80",x"80",x"9C",x"C2",x"47",x"85",x"0C",x"98",x"48",x"96",x"9C",x"7B",x"EE",x"04",x"4B",x"19",x"2E",x"BA",x"14",x"9E",x"D3",x"4F",x"DA",x"FB",x"B9",x"A4",x"30",x"21",x"1C",x"72",x"00",x"79",x"D3",x"B5",x"04",x"38",x"6E",x"7E",x"0F",x"0E",x"40",x"1B",x"1F",x"68",x"9C",x"EF",x"01",x"3C",x"41",x"3F",x"70",x"00",x"C5",x"6E",x"F2",x"FD",x"24",x"0F",x"98",x"3C",x"54",x"53",x"E4",x"17",x"88",x"19",x"13",x"19",x"32",x"C6",x"68",x"A5",x"2C",x"CC",x"AF",x"0A",x"3E",x"E1",x"10",x"96",x"81",x"0A",x"36",x"29",x"9B",x"32",x"B9",x"67",x"99",x"6E",x"B2",x"10",x"D8",x"C9",x"37",x"00",x"3D",x"07",x"B9",x"A9",x"D1",x"B2",x"58",x"06",x"B1",x"83",x"E3",x"27",x"21",x"B2",x"55",x"D3",x"22",x"DE",x"43",x"54",x"C4",x"00",x"E4",x"39",x"86",x"E5",x"E5",x"45",x"12",x"D3",x"70",x"13",x"80",x"B7",x"DB",x"2C",x"9D",x"C0",x"5D",x"86",x"21",x"A1",x"38",x"66",x"51",x"4E",x"C4",x"6F",x"54",x"0E",x"99",x"B8",x"5C",x"89",x"FD",x"04",x"B2",x"72",x"D0",x"D6",x"35",x"D5",x"00",x"76",x"AD",x"21",x"7A",x"E0",x"13",x"43",x"CB",x"7C",x"72",x"66",x"B5",x"C0",x"1A",x"F4",x"83",x"00",x"25",x"A9",x"AB",x"24",x"91",x"D4",x"D5",x"23",x"48",x"AD",x"22",x"7A",x"E9",x"AF",x"69",x"21",x"14",x"86",x"01",x"9F",x"18",x"98",x"DE",x"53",x"0E",x"1F",x"B9",x"EE",x"D0",x"AA",x"8F",x"10",x"43",x"7B",x"1D",x"22",x"32",x"1C",x"9E",x"D5",x"D0",x"80",x"05",x"AA",x"6F",x"AF",x"85",x"4F",x"ED",x"9D",x"71",x"1E",x"ED",x"BE",x"41",x"4D",x"40",x"03",x"56",x"0C",x"75",x"71",x"5B",x"F1",x"04",x"C7",x"50",x"D4",x"8D",x"2D",x"9D",x"F5",x"10",x"C3",x"A8",x"A0",x"8C",x"AA",x"98",x"A0",x"24",x"4D",x"FC",x"65",x"31",x"5B",x"7A",x"00",x"31",x"A9",x"55",x"C6",x"FC",x"B7",x"28",x"E1",x"1D",x"7B",x"03",x"27",x"AE",x"AF",x"B4",x"D8",x"C6",x"4F",x"38",x"94",x"16",x"4D",x"52",x"12",x"4F",x"48",x"23",x"39",x"69",x"8A",x"7A",x"44",x"14",x"C2",x"2F",x"E5",x"F4",x"98",x"B8",x"4F",x"42",x"37",x"CA",x"09",x"30",x"24",x"DA",x"C4",x"3A",x"96",x"7B",x"03",x"2B",x"04",x"E5",x"5E",x"CD",x"4F",x"C5",x"8F",x"AD",x"73",x"A7",x"25",x"13",x"39",x"09",x"06",x"BC",x"A0",x"7D",x"67",x"B9",x"15",x"7D",x"29",x"10",x"7C",x"92",x"02",x"21",x"7B",x"AD",x"A5",x"7A",x"77",x"67",x"BB",x"AC",x"4D",x"B6",x"A6",x"B2",x"B1",x"9E",x"B0",x"A7",x"D6",x"AF",x"79",x"22",x"46",x"54",x"A9",x"55",x"F7",x"56",x"3C",x"10",x"99",x"5F",x"B6",x"A5",x"22",x"B5",x"91",x"54",x"24",x"B4",x"52",x"2E",x"72",x"79",x"5B",x"58",x"59",x"EF",x"5A",x"59",x"89",x"23",x"E6",x"31",x"72",x"F4",x"45",x"83",x"54",x"23",x"97",x"05",x"48",x"4C",x"3B",x"88",x"60",x"95",x"89",x"C4",x"E3",x"ED",x"07",x"48",x"29",x"01",x"CD",x"6B",x"39",x"71",x"9E",x"17",x"4C",x"42",x"6A",x"CF",x"E6",x"42",x"11",x"78",x"5C",x"20",x"9F",x"99",x"60",x"7D",x"9F",x"4D",x"2D",x"E9",x"C5",x"A1",x"9C",x"6B",x"7D",x"88",x"F7",x"DB",x"23",x"42",x"24",x"F0",x"CF",x"20",x"7F",x"B9",x"0D",x"E7",x"C9",x"C0",x"3B",x"06",x"59",x"AA",x"A5",x"80",x"30",x"DC",x"D3",x"A2",x"52",x"3A",x"AB",x"49",x"BD",x"A2",x"00",x"C8",x"44",x"F0",x"F5",x"54",x"63",x"DD",x"80",x"9A",x"20",x"39",x"DE",x"11",x"08",x"9B",x"DF",x"C5",x"86",x"0D",x"E8",x"25",x"B7",x"79",x"D9",x"DD",x"73",x"FC",x"05",x"87",x"98",x"57",x"40",x"77",x"50",x"6B",x"E6",x"E6",x"28",x"69",x"41",x"55",x"0E",x"B4",x"FD",x"56",x"60",x"6A",x"0C",x"18",x"15",x"37",x"62",x"76",x"50",x"08",x"2B",x"A7",x"E0",x"A6",x"79",x"A5",x"A4",x"5E",x"99",x"DC",x"B1",x"C8",x"73",x"6E",x"01",x"9B",x"B3",x"B4",x"05",x"81",x"C8",x"0D",x"64",x"25",x"0A",x"41",x"5C",x"D7",x"5D",x"7B",x"5E",x"CE",x"6C",x"84",x"C5",x"DC",x"5E",x"15",x"76",x"0D",x"6B",x"99",x"0E",x"6C",x"25",x"90",x"65",x"70",x"B1",x"D9",x"1E",x"A0",x"1F",x"5B",x"D4",x"5A",x"F3",x"59",x"58",x"BC",x"53",x"7F",x"68",x"F0",x"54",x"A5",x"FB",x"F0",x"46",x"53",x"3D",x"52",x"51",x"CF",x"AA",x"E9",x"01",x"1C",x"FA",x"1C",x"4F",x"E1",x"5F",x"7A",x"5E",x"5D",x"9E",x"89",x"AB",x"90",x"56",x"66",x"3D",x"5C",x"5A",x"7D",x"82",x"56",x"91",x"63",x"66",x"26",x"B6",x"52",x"02",x"30",x"61",x"6C",x"C6",x"C4",x"91",x"82",x"46",x"BE",x"01",x"64",x"80",x"11",x"F9",x"5C",x"5A",x"73",x"3A",x"2B",x"41",x"57",x"3D",x"56",x"37",x"65",x"55",x"53",x"AD",x"54",x"5A",x"8D",x"50",x"5A",x"8E",x"51",x"FA",x"52",x"14",x"94",x"53",x"7D",x"7D",x"67",x"F6",x"C6",x"5B",x"22",x"3C",x"F4",x"39",x"AF",x"62",x"71",x"C9",x"E5",x"56",x"B9",x"2E",x"95",x"E3",x"D9",x"B5",x"99",x"4A",x"59",x"CE",x"50",x"78",x"28",x"57",x"6B",x"08",x"CA",x"0C",x"E1",x"C8",x"3C",x"00",x"5C",x"CD",x"18",x"02",x"01",x"30",x"28",x"83",x"84",x"8A",x"32",x"2C",x"1C",x"91",x"BE",x"44",x"DC",x"D0",x"BD",x"4F",x"99",x"59",x"72",x"02",x"9A",x"CF",x"4A",x"1F",x"20",x"A0",x"49",x"8D",x"F8",x"D7",x"8E",x"A5",x"D8",x"04",x"6F",x"D9",x"A5",x"04",x"62",x"DA",x"32",x"6E",x"E0",x"50",x"03",x"57",x"C9",x"09",x"B2",x"B0",x"B0",x"14",x"EC",x"B0",x"ED",x"28",x"C0",x"0F",x"C0",x"0A",x"6F",x"64",x"80",x"11",x"99",x"66",x"16",x"E1",x"06",x"31",x"69",x"0A",x"F7",x"13",x"58",x"81",x"0A",x"60",x"74",x"A5",x"EB",x"20",x"6E",x"C0",x"52",x"21",x"E1",x"C9",x"5A",x"1C",x"B2",x"F5",x"25",x"08",x"B3",x"02",x"30",x"B1",x"0E",x"54",x"D4",x"2D",x"F0",x"E1",x"D3",x"B6",x"AE",x"31",x"2C",x"D9",x"9D",x"C9",x"72",x"DB",x"01",x"55",x"AE",x"25",x"A6",x"46",x"ED",x"5D",x"55",x"A4",x"52",x"59",x"E1",x"0F",x"46",x"E7",x"FA",x"73",x"C1",x"09",x"03",x"46",x"A6",x"03",x"04",x"6C",x"6E",x"38",x"73",x"90",x"F2",x"80",x"7D",x"E8",x"45",x"16",x"B0",x"2F",x"00",x"F0",x"71",x"AA",x"1D",x"1C",x"20",x"FB",x"16",x"F3",x"80",x"07",x"EC",x"23",x"4C",x"EA",x"FD",x"0A",x"13",x"03",x"F0",x"86",x"9F",x"F1",x"9E",x"D4",x"30",x"9D",x"A5",x"9C",x"5A",x"B5",x"4E",x"26",x"16",x"60",x"A8",x"E3",x"A9",x"6D",x"19",x"A3",x"49",x"29",x"C0",x"48",x"44",x"33",x"A3",x"AE",x"A1",x"78",x"CB",x"77",x"B5",x"06",x"9C",x"99",x"3B",x"82",x"07",x"B3",x"E6",x"0B",x"9C",x"EB",x"66",x"9E",x"01",x"E8",x"EB",x"82",x"C7",x"D1",x"27",x"BA",x"05",x"8D",x"1E",x"EC",x"06",x"F3",x"D3",x"04",x"D8",x"64",x"70",x"03",x"A1",x"87",x"6A",x"B0",x"8D",x"0A",x"7A",x"00",x"7E",x"DD",x"11",x"05",x"68",x"A9",x"8A",x"C8",x"58",x"70",x"BD",x"32",x"EE",x"AC",x"36",x"B4",x"3F",x"95",x"20",x"BC",x"3C",x"40",x"13",x"7C",x"8D",x"68",x"07",x"2F",x"6A",x"11",x"FC",x"CA",x"A5",x"AD",x"E6",x"96",x"76",x"37",x"9A",x"2A",x"CB",x"4B",x"B5",x"6D",x"02",x"CE",x"A0",x"B1",x"22",x"75",x"A5",x"6E",x"99",x"A7",x"D0",x"AA",x"F7",x"47",x"00",x"8C",x"79",x"BD",x"2E",x"06",x"59",x"F1",x"8B",x"0D",x"BA",x"E8",x"5A",x"73",x"2B",x"18",x"0F",x"74",x"56",x"D2",x"6A",x"D6",x"32",x"83",x"41",x"50",x"CC",x"71",x"6B",x"02",x"42",x"40",x"E3",x"41",x"7F",x"BC",x"8B",x"C9",x"4F",x"20",x"59",x"34",x"F1",x"D5",x"54",x"16",x"01",x"42",x"D9",x"02",x"A7",x"4A",x"19",x"FF",x"AD",x"7C",x"35",x"07",x"21",x"D8",x"44",x"2E",x"C2",x"74",x"53",x"B9",x"18",x"70",x"0C",x"AC",x"6B",x"B7",x"DE",x"DD",x"9E",x"DC",x"E7",x"DB",x"08",x"BD",x"E2",x"E7",x"E1",x"C9",x"61",x"E0",x"4A",x"DF",x"B5",x"65",x"45",x"53",x"27",x"BC",x"9B",x"6A",x"C0",x"EA",x"A4",x"E9",x"EB",x"E7",x"DB",x"E8",x"94",x"AD",x"E7",x"7C",x"FE",x"AA",x"14",x"7D",x"FA",x"6D",x"40",x"BC",x"85",x"85",x"1E",x"35",x"AD",x"D3",x"73",x"D9",x"FA",x"7E",x"FE",x"D4",x"46",x"84",x"2C",x"87",x"4A",x"62",x"D7",x"F0",x"0A",x"63",x"4C",x"7E",x"77",x"BE",x"64",x"56",x"26",x"9B",x"1C",x"41",x"2F",x"60",x"CE",x"80",x"04",x"AA",x"DD",x"0F",x"C8",x"B9",x"BC",x"F5",x"73",x"D9",x"BB",x"7C",x"F0",x"F4",x"3E",x"01",x"B0",x"02",x"9D",x"D2",x"B1",x"A9",x"47",x"13",x"B4",x"F0",x"70",x"D6",x"01",x"57",x"73",x"5D",x"C3",x"D4",x"08",x"34",x"72",x"05",x"25",x"80",x"06",x"C8",x"08",x"D5",x"4C",x"F3",x"29",x"EF",x"20",x"40",x"08",x"0E",x"9F",x"4F",x"07",x"AF",x"96",x"27",x"B4",x"25",x"4C",x"FC",x"63",x"7E",x"47",x"25",x"53",x"8D",x"CC",x"2F",x"D0",x"75",x"87",x"2F",x"F6",x"46",x"55",x"61",x"36",x"A4",x"31",x"40",x"AA",x"6A",x"B4",x"3A",x"84",x"66",x"B6",x"F1",x"03",x"2B",x"6B",x"21",x"77",x"79",x"9E",x"9E",x"78",x"4C",x"A9",x"79",x"45",x"D3",x"54",x"B1",x"A9",x"9B",x"2D",x"AC",x"A7",x"04",x"C0",x"B7",x"18",x"90",x"17",x"7E",x"A9",x"D6",x"AE",x"F8",x"E2",x"32",x"74",x"89",x"49",x"76",x"B5",x"CE",x"7E",x"5A",x"6F",x"04",x"CA",x"99",x"19",x"A0",x"AC",x"57",x"10",x"9B",x"21",x"C0",x"43",x"B6",x"43",x"E2",x"48",x"0E",x"DC",x"A9",x"BB",x"81",x"9D",x"36",x"2C",x"A7",x"31",x"A0",x"72",x"4E",x"8D",x"80",x"DD",x"6D",x"CC",x"75",x"43",x"47",x"76",x"3B",x"31",x"96",x"0C",x"DB",x"48",x"7B",x"09",x"A0",x"25",x"09",x"77",x"B8",x"31",x"0B",x"05",x"5C",x"0F",x"3C",x"05",x"1F",x"05",x"A8",x"30",x"07",x"74",x"B8",x"8F",x"0B",x"5A",x"6C",x"A9",x"4E",x"57",x"6D",x"AD",x"6E",x"EC",x"1A",x"8D",x"6F",x"F4",x"9F",x"F0",x"C1",x"02",x"70",x"F5",x"71",x"B0",x"A9",x"03",x"D4",x"72",x"95",x"64",x"7B",x"59",x"74",x"89",x"DA",x"69",x"73",x"56",x"05",x"FB",x"75",x"4D",x"9C",x"76",x"E9",x"93",x"FF",x"8A",x"C2",x"20",x"8F",x"64",x"8D",x"78",x"3F",x"A4",x"79",x"9D",x"50",x"A5",x"F0",x"54",x"8D",x"93",x"B6",x"25",x"D0",x"6C",x"69",x"24",x"1A",x"59",x"AA",x"BC",x"47",x"19",x"E0",x"79",x"56",x"BC",x"65",x"A8",x"F0",x"89",x"AB",x"0C",x"7A",x"7D",x"5C",x"D6",x"2E",x"4C",x"10",x"64",x"3D",x"48",x"51",x"02",x"9C",x"A5",x"04",x"F9",x"A9",x"8E",x"01",x"DF",x"A9",x"6C",x"D4",x"8D",x"05",x"D7",x"67",x"99",x"72",x"58",x"DC",x"71",x"97",x"E0",x"5A",x"31",x"61",x"7B",x"18",x"D0",x"AD",x"76",x"66",x"C3",x"29",x"FC",x"2E",x"01",x"27",x"00",x"48",x"AD",x"51",x"64",x"C3",x"09",x"03",x"8E",x"AD",x"02",x"DD",x"9C",x"20",x"F5",x"06",x"B7",x"21",x"52",x"2D",x"8D",x"16",x"D0",x"EA",x"28",x"0A",x"03",x"50",x"EB",x"51",x"32",x"2C",x"94",x"42",x"B6",x"B3",x"2D",x"D0",x"6C",x"5C",x"AD",x"12",x"47",x"51",x"35",x"07",x"CA",x"D0",x"AA",x"37",x"01",x"CB",x"CC",x"94",x"AE",x"CD",x"55",x"BE",x"33",x"39",x"4B",x"00",x"71",x"88",x"02",x"61",x"45",x"08",x"01",x"4C",x"27",x"B1",x"E8",x"08",x"9C",x"9A",x"CF",x"8E",x"A5",x"D0",x"A9",x"1F",x"D1",x"92",x"FA",x"21",x"D2",x"9C",x"A5",x"D3",x"78",x"B1",x"C7",x"82",x"56",x"3D",x"21",x"4F",x"2A",x"2B",x"9E",x"D4",x"DA",x"8A",x"77",x"06",x"FC",x"71",x"69",x"B2",x"0A",x"DE",x"ED",x"9C",x"8B",x"D2",x"8D",x"DE",x"F3",x"7D",x"8A",x"87",x"A1",x"8E",x"9B",x"8D",x"F1",x"E7",x"BB",x"8C",x"29",x"AD",x"8B",x"7D",x"03",x"9D",x"12",x"92",x"97",x"44",x"B9",x"F0",x"3B",x"AA",x"94",x"5A",x"80",x"B0",x"42",x"EA",x"50",x"20",x"E2",x"85",x"AC",x"6F",x"32",x"5C",x"DF",x"26",x"E5",x"8B",x"A1",x"06",x"26",x"8A",x"B4",x"63",x"C9",x"4F",x"D4",x"02",x"4A",x"BF",x"D3",x"42",x"C8",x"9C",x"09",x"76",x"B1",x"05",x"D9",x"48",x"0F",x"DB",x"B1",x"30",x"CE",x"A2",x"61",x"A5",x"8D",x"44",x"CA",x"AF",x"C2",x"9F",x"C0",x"51",x"A5",x"80",x"AF",x"05",x"02",x"D6",x"18",x"44",x"A6",x"96",x"10",x"29",x"C9",x"79",x"2D",x"7A",x"24",x"98",x"20",x"03",x"E0",x"89",x"A5",x"04",x"E1",x"05",x"04",x"E2",x"1C",x"37",x"DE",x"0B",x"DA",x"98",x"49",x"88",x"84",x"05",x"ED",x"8B",x"10",x"D0",x"52",x"39",x"C5",x"C8",x"8F",x"05",x"06",x"A2",x"1C",x"00",x"15",x"A8",x"75",x"07",x"90",x"FB",x"24",x"60",x"7E",x"B7",x"88",x"26",x"28",x"62",x"C6",x"23",x"E2",x"07",x"FA",x"1A",x"B8",x"23",x"9A",x"E9",x"E7",x"8C",x"38",x"D9",x"61",x"66",x"C2",x"A3",x"0E",x"5C",x"D4",x"25",x"61",x"EF",x"2E",x"F1",x"30",x"48",x"0D",x"AC",x"DD",x"C7",x"48",x"4E",x"2A",x"29",x"6B",x"EC",x"9C",x"96",x"85",x"6E",x"69",x"10",x"B0",x"74",x"7F",x"4A",x"29",x"01",x"F0",x"5A",x"9C",x"7E",x"DC",x"A9",x"04",x"8D",x"FE",x"54",x"80",x"B0",x"4B",x"71",x"AF",x"0A",x"7F",x"0A",x"17",x"8B",x"E3",x"20",x"36",x"8E",x"DA",x"6E",x"6E",x"F8",x"88",x"3D",x"A2",x"66",x"C9",x"93",x"65",x"04",x"4E",x"9C",x"69",x"CE",x"F4",x"F2",x"46",x"90",x"0B",x"65",x"0C",x"23",x"81",x"85",x"52",x"CE",x"56",x"87",x"49",x"AC",x"51",x"14",x"88",x"B2",x"99",x"DA",x"CE",x"59",x"41",x"AE",x"24",x"6B",x"4A",x"B0",x"4C",x"8A",x"9D",x"0D",x"6A",x"B6",x"89",x"AA",x"9C",x"74",x"85",x"85",x"22",x"1E",x"A9",x"7F",x"A2",x"FC",x"64",x"14",x"09",x"81",x"30",x"89",x"52",x"DB",x"D4",x"61",x"04",x"5C",x"74",x"AC",x"64",x"0A",x"EA",x"22",x"C9",x"0A",x"59",x"E5",x"B7",x"CA",x"75",x"80",x"8B",x"21",x"2B",x"81",x"15",x"ED",x"58",x"82",x"A5",x"E0",x"8D",x"83",x"DE",x"52",x"CC",x"D0",x"9C",x"2C",x"19",x"EE",x"C9",x"05",x"D9",x"B0",x"20",x"80",x"DB",x"18",x"6D",x"E3",x"64",x"96",x"95",x"AC",x"F1",x"B9",x"7F",x"D8",x"92",x"0A",x"D4",x"86",x"35",x"A4",x"D9",x"00",x"C5",x"A7",x"E2",x"16",x"78",x"89",x"25",x"12",x"40",x"58",x"AD",x"3D",x"D2",x"05",x"92",x"08",x"95",x"29",x"14",x"1F",x"8E",x"55",x"17",x"12",x"08",x"ED",x"D3",x"95",x"50",x"1B",x"48",x"AC",x"CE",x"4D",x"99",x"2E",x"FA",x"67",x"80",x"07",x"BB",x"4C",x"72",x"49",x"8A",x"08",x"4D",x"5C",x"30",x"A8",x"B8",x"AC",x"4C",x"E7",x"93",x"8E",x"3C",x"93",x"66",x"C9",x"0D",x"35",x"C6",x"D0",x"0B",x"0D",x"0D",x"FC",x"C4",x"A5",x"63",x"26",x"08",x"F0",x"91",x"F0",x"B9",x"1F",x"41",x"64",x"C2",x"41",x"93",x"00",x"07",x"1F",x"A3",x"F5",x"69",x"65",x"0F",x"62",x"05",x"94",x"34",x"5C",x"C7",x"0D",x"33",x"0A",x"80",x"83",x"32",x"D0",x"48",x"84",x"49",x"80",x"31",x"B6",x"9A",x"07",x"C2",x"4C",x"04",x"12",x"6E",x"63",x"2C",x"1D",x"6C",x"2B",x"03",x"0D",x"21",x"F8",x"59",x"66",x"98",x"72",x"A2",x"07",x"C8",x"C9",x"38",x"C8",x"05",x"45",x"87",x"21",x"54",x"45",x"BF",x"50",x"B1",x"50",x"08",x"30",x"8B",x"46",x"D5",x"1A",x"41",x"4C",x"9B",x"05",x"3B",x"5F",x"15",x"A0",x"EB",x"B0",x"D5",x"C1",x"41",x"9C",x"38",x"4A",x"EE",x"A8",x"08",x"F7",x"19",x"7E",x"27",x"D0",x"F6",x"A1",x"84",x"06",x"50",x"9A",x"C9",x"23",x"6E",x"D8",x"54",x"43",x"49",x"80",x"03",x"9C",x"B9",x"B0",x"83",x"F8",x"D4",x"BB",x"5F",x"44",x"5D",x"4D",x"66",x"C2",x"2F",x"1B",x"04",x"80",x"06",x"A2",x"08",x"DE",x"D5",x"01",x"4A",x"69",x"98",x"2E",x"01",x"D3",x"82",x"2D",x"37",x"C9",x"14",x"F0",x"F8",x"C7",x"4D",x"36",x"AE",x"F2",x"CB",x"EA",x"1C",x"79",x"E5",x"E3",x"03",x"E6",x"00",x"89",x"9F",x"51",x"A9",x"80",x"50",x"D0",x"F0",x"00",x"18",x"AD",x"67",x"99",x"7B",x"88",x"32",x"4A",x"0C",x"28",x"37",x"6C",x"C9",x"0D",x"D0",x"EC",x"C8",x"A3",x"1D",x"3B",x"86",x"A0",x"4C",x"39",x"37",x"73",x"1A",x"02",x"93",x"BA",x"66",x"3E",x"7C",x"6E",x"E1",x"95",x"01",x"C8",x"02",x"60",x"5B",x"06",x"ED",x"6C",x"1B",x"2C",x"14",x"E0",x"07",x"AA",x"6B",x"D2",x"16",x"F8",x"8C",x"75",x"23",x"DB",x"3A",x"8E",x"05",x"12",x"C2",x"A2",x"80",x"C5",x"A7",x"49",x"DC",x"66",x"76",x"A7",x"38",x"F8",x"E4",x"9A",x"E8",x"04",x"67",x"9C",x"09",x"E6",x"E8",x"35",x"A7",x"6D",x"C8",x"C0",x"CE",x"2C",x"C7",x"10",x"D6",x"EF",x"65",x"CD",x"6C",x"8F",x"E6",x"76",x"34",x"A0",x"F7",x"E9",x"60",x"53",x"0B",x"61",x"73",x"58",x"E3",x"62",x"23",x"E5",x"0B",x"08",x"3D",x"C2",x"68",x"76",x"7B",x"0A",x"08",x"B2",x"05",x"B4",x"1E",x"06",x"04",x"99",x"0C",x"1B",x"E3",x"79",x"61",x"6C",x"5A",x"D1",x"95",x"D9",x"11",x"52",x"F1",x"5D",x"81",x"B8",x"38",x"9D",x"0B",x"F1",x"8E",x"24",x"80",x"4D",x"43",x"E7",x"AC",x"6D",x"07",x"43",x"97",x"4E",x"2E",x"18",x"CD",x"0C",x"5F",x"94",x"E1",x"A7",x"4E",x"C8",x"15",x"CD",x"87",x"15",x"6B",x"36",x"0B",x"3C",x"C5",x"1F",x"07",x"27",x"93",x"C3",x"A9",x"8F",x"F1",x"3E",x"15",x"90",x"1C",x"99",x"D0",x"AD",x"05",x"70",x"35",x"D1",x"B0",x"A9",x"37",x"88",x"10",x"9F",x"D9",x"EA",x"65",x"42",x"2C",x"32",x"F2",x"04",x"48",x"5C",x"6A",x"0E",x"6D",x"CA",x"20",x"87",x"2D",x"2C",x"0A",x"3E",x"57",x"59",x"C2",x"B1",x"12",x"B6",x"DE",x"34",x"22",x"1B",x"96",x"2F",x"9C",x"2B",x"4B",x"21",x"F0",x"27",x"70",x"8E",x"EA",x"21",x"1E",x"9C",x"E3",x"42",x"1E",x"E4",x"F0",x"89",x"87",x"42",x"80",x"C6",x"AE",x"8E",x"BD",x"3A",x"99",x"6E",x"91",x"EE",x"1E",x"A2",x"87",x"BB",x"AC",x"9E",x"8F",x"BD",x"7D",x"CE",x"53",x"F4",x"CA",x"0B",x"F8",x"66",x"01",x"8A",x"80",x"24",x"FF",x"90",x"10",x"01",x"E6",x"80",x"3A",x"59",x"6C",x"22",x"9B",x"A1",x"21",x"8D",x"50",x"EF",x"9C",x"80",x"FE",x"E5",x"90",x"86",x"37",x"8D",x"5B",x"31",x"30",x"7A",x"75",x"B6",x"A4",x"4D",x"D9",x"C2",x"75",x"2D",x"AD",x"93",x"4E",x"79",x"27",x"2B",x"5C",x"5D",x"A5",x"A9",x"92",x"26",x"2C",x"A7",x"E6",x"EA",x"09",x"2A",x"63",x"AE",x"80",x"19",x"83",x"1C",x"80",x"A4",x"03",x"8D",x"43",x"D6",x"18",x"7F",x"CB",x"98",x"A0",x"52",x"B1",x"5C",x"E1",x"0A",x"D0",x"D9",x"23",x"75",x"1C",x"78",x"D7",x"35",x"0F",x"92",x"CA",x"39",x"7C",x"32",x"E4",x"60",x"30",x"52",x"31",x"08",x"35",x"41",x"A3",x"2F",x"36",x"CB",x"D4",x"0E",x"80",x"40",x"FF",x"A7",x"B7",x"81",x"2E",x"18",x"A0",x"06",x"4E",x"48",x"8A",x"64",x"EC",x"34",x"F1",x"B2",x"83",x"B1",x"42",x"5B",x"39",x"5D",x"3E",x"82",x"C5",x"25",x"CB",x"22",x"EE",x"5A",x"51",x"3E",x"81",x"11",x"88",x"C6",x"63",x"BE",x"3E",x"C5",x"2C",x"BC",x"AE",x"90",x"63",x"79",x"89",x"7D",x"23",x"FA",x"8D",x"CB",x"1F",x"C9",x"59",x"CA",x"5C",x"B9",x"7F",x"39",x"5C",x"0D",x"98",x"2B",x"F5",x"8D",x"B8",x"99",x"25",x"9A",x"A7",x"84",x"BF",x"06",x"A5",x"7A",x"A9",x"01",x"F6",x"86",x"80",x"1B",x"DC",x"9B",x"08",x"71",x"38",x"F3",x"B3",x"03",x"AF",x"8D",x"55",x"66",x"21",x"9C",x"95",x"DD",x"CD",x"D8",x"9D",x"59",x"D0",x"D8",x"DB",x"9B",x"90",x"47",x"AE",x"F0",x"89",x"69",x"9C",x"F9",x"80",x"B1",x"10",x"A9",x"0A",x"EF",x"30",x"8C",x"7D",x"6D",x"10",x"25",x"D9",x"29",x"F0",x"D0",x"EA",x"F3",x"49",x"49",x"6D",x"0A",x"8D",x"96",x"C7",x"D8",x"9E",x"95",x"7D",x"6A",x"C9",x"BE",x"25",x"2F",x"C7",x"5D",x"08",x"6C",x"2A",x"1C",x"92",x"CE",x"28",x"01",x"C8",x"AC",x"A2",x"90",x"43",x"88",x"36",x"03",x"BC",x"60",x"04",x"50",x"C3",x"97",x"C0",x"FD",x"34",x"07",x"F8",x"4C",x"AC",x"17",x"C2",x"C1",x"95",x"F2",x"52",x"36",x"09",x"11",x"40",x"C0",x"2B",x"DD",x"02",x"B5",x"0E",x"4E",x"F0",x"0A",x"D5",x"C9",x"21",x"46",x"A3",x"54",x"3C",x"7C",x"BA",x"01",x"71",x"1A",x"D8",x"00",x"98",x"11",x"C0",x"10",x"39",x"01",x"13",x"12",x"78",x"96",x"40",x"35",x"B8",x"38",x"0D",x"80",x"14",x"EB",x"0A",x"3F",x"81",x"80",x"3C",x"88",x"DF",x"03",x"18",x"34",x"C8",x"37",x"44",x"F0",x"1A",x"3A",x"04",x"01",x"3A",x"0C",x"B1",x"AD",x"2F",x"44",x"6C",x"26",x"53",x"7F",x"0D",x"B0",x"1F",x"4D",x"1F",x"02",x"33",x"13",x"81",x"24",x"BE",x"85",x"95",x"03",x"1A",x"82",x"14",x"C0",x"04",x"C6",x"40",x"08",x"15",x"3C",x"29",x"64",x"EE",x"E3",x"04",x"61",x"80",x"64",x"16",x"83",x"21",x"42",x"3C",x"3A",x"AD",x"38",x"10",x"20",x"B5",x"69",x"A2",x"71",x"F9",x"FD",x"75",x"27",x"92",x"15",x"17",x"FF",x"A7",x"39",x"29",x"4B",x"41",x"5F",x"6A",x"C9",x"90",x"E9",x"A5",x"43",x"B9",x"52",x"FA",x"72",x"0B",x"2F",x"20",x"12",x"F0",x"92",x"07",x"2E",x"11",x"0B",x"1E",x"A7",x"08",x"9F",x"F0",x"3D",x"CB",x"94",x"EC",x"E0",x"02",x"AB",x"33",x"DD",x"C5",x"05",x"3B",x"23",x"44",x"7B",x"9C",x"01",x"11",x"02",x"E2",x"66",x"5F",x"BF",x"8B",x"D0",x"86",x"F6",x"80",x"B6",x"B1",x"87",x"C7",x"54",x"B0",x"63",x"C6",x"4F",x"69",x"D0",x"45",x"87",x"E0",x"54",x"00",x"08",x"2A",x"34",x"99",x"0A",x"D0",x"11",x"36",x"38",x"09",x"70",x"37",x"05",x"F1",x"1A",x"AC",x"80",x"94",x"65",x"DA",x"C8",x"E8",x"12",x"3E",x"71",x"B3",x"04",x"05",x"84",x"61",x"50",x"82",x"4F",x"1C",x"34",x"50",x"E0",x"54",x"43",x"7B",x"6C",x"E0",x"C2",x"64",x"07",x"25",x"05",x"B3",x"F5",x"B2",x"3C",x"B1",x"0B",x"B0",x"78",x"DD",x"09",x"AD",x"27",x"5C",x"EA",x"C0",x"80",x"15",x"B9",x"A2",x"98",x"C8",x"38",x"7A",x"BD",x"3C",x"89",x"B3",x"35",x"44",x"DA",x"76",x"47",x"16",x"9C",x"69",x"79",x"26",x"76",x"0B",x"A1",x"E9",x"CF",x"C1",x"4E",x"B9",x"99",x"87",x"B4",x"E4",x"AC",x"28",x"AB",x"AA",x"CF",x"A9",x"53",x"A8",x"B6",x"78",x"5B",x"6F",x"8A",x"3F",x"31",x"EF",x"1A",x"44",x"40",x"7B",x"84",x"57",x"70",x"5A",x"48",x"9A",x"6A",x"B0",x"08",x"03",x"AB",x"3F",x"B5",x"1F",x"15",x"44",x"9D",x"C1",x"01",x"C6",x"0E",x"02",x"38",x"52",x"FF",x"00",x"7C",x"0F",x"91",x"03",x"1E",x"E4",x"15",x"B0",x"1D",x"5A",x"4A",x"69",x"0D",x"23",x"21",x"35",x"E8",x"B3",x"08",x"07",x"4F",x"CE",x"C5",x"C5",x"A4",x"E5",x"6E",x"27",x"0E",x"D5",x"7E",x"C6",x"6C",x"B5",x"AF",x"3E",x"70",x"ED",x"3A",x"A8",x"2B",x"65",x"A4",x"EC",x"0F",x"4A",x"09",x"76",x"8F",x"0E",x"A8",x"16",x"14",x"1A",x"F1",x"6F",x"5C",x"77",x"5B",x"3E",x"0B",x"AE",x"2C",x"45",x"08",x"95",x"91",x"D7",x"9F",x"77",x"95",x"71",x"94",x"42",x"80",x"57",x"9F",x"34",x"1A",x"05",x"BF",x"62",x"3D",x"50",x"17",x"2C",x"61",x"14",x"F1",x"B9",x"75",x"D9",x"55",x"B4",x"61",x"B3",x"76",x"4B",x"E6",x"A5",x"34",x"E5",x"48",x"4A",x"83",x"E4",x"94",x"E3",x"AA",x"7C",x"BF",x"67",x"AF",x"02",x"CE",x"33",x"02",x"CD",x"13",x"49",x"AD",x"AC",x"78",x"3F",x"47",x"29",x"03",x"FC",x"68",x"9E",x"44",x"3A",x"38",x"1C",x"06",x"C8",x"41",x"84",x"1A",x"D0",x"70",x"07",x"02",x"24",x"21",x"30",x"00",x"19",x"F6",x"DF",x"3B",x"B2",x"21",x"22",x"03",x"92",x"C1",x"48",x"C0",x"3C",x"0A",x"05",x"79",x"48",x"68",x"D0",x"04",x"1A",x"FA",x"03",x"8A",x"38",x"F2",x"5D",x"4F",x"DE",x"05",x"69",x"CF",x"FA",x"9A",x"99",x"2C",x"3E",x"BD",x"62",x"99",x"AF",x"90",x"85",x"3A",x"B4",x"01",x"14",x"D6",x"83",x"92",x"11",x"9C",x"19",x"B5",x"F0",x"2F",x"B8",x"09",x"36",x"07",x"E0",x"56",x"A9",x"3F",x"BF",x"63",x"44",x"09",x"83",x"8C",x"67",x"6E",x"80",x"0F",x"41",x"32",x"DB",x"2E",x"40",x"C5",x"70",x"88",x"11",x"67",x"F2",x"BB",x"50",x"CC",x"1F",x"59",x"95",x"6E",x"4D",x"C5",x"0B",x"B6",x"80",x"82",x"3B",x"5E",x"4C",x"15",x"CB",x"2B",x"1B",x"91",x"6B",x"89",x"14",x"1C",x"5A",x"26",x"63",x"1B",x"FB",x"31",x"02",x"79",x"38",x"0A",x"8E",x"89",x"B2",x"0C",x"62",x"9B",x"69",x"CF",x"A5",x"48",x"9D",x"4E",x"27",x"AF",x"B9",x"6B",x"75",x"3D",x"77",x"37",x"F8",x"4D",x"2C",x"4D",x"E0",x"CB",x"6B",x"71",x"D4",x"74",x"1C",x"54",x"48",x"E4",x"12",x"4B",x"90",x"09",x"D2",x"8C",x"47",x"C9",x"D9",x"D0",x"E2",x"44",x"5C",x"E2",x"44",x"6A",x"D6",x"A0",x"34",x"24",x"61",x"91",x"CE",x"43",x"31",x"9C",x"26",x"00",x"60",x"CE",x"F3",x"FD",x"48",x"BF",x"43",x"C2",x"76",x"19",x"08",x"B0",x"30",x"57",x"64",x"8F",x"40",x"17",x"B5",x"60",x"56",x"CC",x"3A",x"ED",x"94",x"80",x"98",x"CA",x"81",x"A9",x"08",x"0F",x"9B",x"98",x"07",x"80",x"19",x"A2",x"99",x"A8",x"B2",x"4C",x"2E",x"9D",x"0A",x"9E",x"3D",x"56",x"6D",x"0D",x"6A",x"03",x"B0",x"4B",x"4C",x"05",x"44",x"08",x"E7",x"40",x"B7",x"3A",x"D4",x"FB",x"8B",x"65",x"03",x"CA",x"EB",x"EE",x"61",x"93",x"08",x"8C",x"8E",x"CF",x"0C",x"8A",x"65",x"73",x"58",x"C5",x"67",x"C8",x"32",x"E9",x"D0",x"E3",x"B0",x"22",x"03",x"BB",x"39",x"48",x"07",x"72",x"66",x"2D",x"89",x"5A",x"47",x"B7",x"28",x"BA",x"31",x"1D",x"E1",x"87",x"5F",x"DF",x"DD",x"A0",x"98",x"62",x"71",x"80",x"2B",x"6C",x"64",x"50",x"F0",x"CB",x"D2",x"99",x"FB",x"0E",x"78",x"9A",x"54",x"68",x"2A",x"6B",x"EC",x"9C",x"3E",x"D0",x"08",x"AA",x"B7",x"6A",x"00",x"67",x"61",x"E3",x"C2",x"05",x"D0",x"6A",x"B6",x"DC",x"03",x"35",x"A8",x"4E",x"61",x"99",x"33",x"8D",x"5C",x"28",x"08",x"28",x"AF",x"7A",x"67",x"D7",x"71",x"5B",x"D5",x"2C",x"8E",x"61",x"39",x"6B",x"09",x"80",x"0C",x"CC",x"46",x"02",x"CC",x"42",x"E6",x"D3",x"82",x"7F",x"80",x"63",x"50",x"C9",x"9C",x"A4",x"CA",x"61",x"39",x"8B",x"0B",x"13",x"DB",x"44",x"47",x"10",x"46",x"95",x"02",x"57",x"61",x"CD",x"A1",x"47",x"66",x"96",x"B0",x"80",x"44",x"49",x"2B",x"C5",x"A6",x"3C",x"5C",x"4A",x"1F",x"C9",x"CD",x"91",x"73",x"CC",x"32",x"14",x"F6",x"A5",x"90",x"DD",x"C0",x"4A",x"9B",x"49",x"78",x"A9",x"51",x"D8",x"20",x"C9",x"62",x"47",x"7C",x"4E",x"00",x"BA",x"BB",x"9B",x"B9",x"CD",x"76",x"6A",x"B0",x"38",x"27",x"51",x"72",x"AC",x"84",x"66",x"CF",x"AD",x"B8",x"78",x"5E",x"A6",x"12",x"D1",x"67",x"11",x"D3",x"F5",x"AD",x"71",x"47",x"82",x"52",x"63",x"9B",x"51",x"C1",x"71",x"02",x"71",x"A3",x"E0",x"90",x"17",x"BA",x"4D",x"01",x"5A",x"06",x"F0",x"5A",x"65",x"C1",x"74",x"B3",x"00",x"55",x"80",x"40",x"C3",x"54",x"F5",x"63",x"5A",x"E4",x"D4",x"F8",x"99",x"4E",x"2A",x"34",x"55",x"C2",x"3E",x"7A",x"5D",x"98",x"1C",x"33",x"4A",x"6A",x"5D",x"F6",x"69",x"0F",x"6F",x"40",x"6B",x"31",x"5C",x"41",x"EE",x"F0",x"B4",x"09",x"9B",x"3A",x"95",x"B4",x"CD",x"93",x"24",x"D3",x"E8",x"20",x"79",x"29",x"7F",x"53",x"EA",x"61",x"D3",x"FC",x"3B",x"6A",x"4E",x"B7",x"5A",x"58",x"C7",x"5B",x"87",x"40",x"63",x"41",x"3C",x"85",x"E3",x"65",x"7F",x"F3",x"51",x"82",x"30",x"60",x"B7",x"E2",x"94",x"E0",x"98",x"F1",x"AE",x"59",x"24",x"46",x"4F",x"AE",x"19",x"C5",x"5C",x"D1",x"EB",x"8A",x"C8",x"F1",x"E9",x"B0",x"3A",x"D5",x"99",x"0E",x"A0",x"5D",x"CC",x"D6",x"17",x"62",x"46",x"4C",x"C7",x"2C",x"67",x"92",x"A4",x"90",x"EB",x"69",x"A6",x"1A",x"64",x"38",x"9E",x"09",x"41",x"51",x"8A",x"F3",x"E9",x"72",x"83",x"40",x"C6",x"5A",x"B0",x"01",x"CA",x"20",x"B3",x"63",x"D0",x"FE",x"23",x"61",x"6B",x"F7",x"AF",x"8E",x"A8",x"29",x"26",x"AA",x"98",x"E0",x"53",x"A2",x"FF",x"86",x"04",x"E5",x"F9",x"59",x"78",x"F8",x"5A",x"8A",x"15",x"A9",x"6A",x"4E",x"AD",x"AF",x"33",x"60",x"6A",x"04",x"69",x"3A",x"7C",x"A9",x"2A",x"50",x"1C",x"2D",x"55",x"6C",x"B0",x"E4",x"01",x"68",x"F5",x"30",x"45",x"A5",x"84",x"8E",x"91",x"5F",x"A4",x"C8",x"44",x"64",x"55",x"AE",x"8A",x"7C",x"58",x"2F",x"54",x"2A",x"4C",x"5A",x"45",x"38",x"AF",x"E2",x"59",x"84",x"C6",x"B5",x"20",x"B2",x"25",x"6E",x"00",x"40",x"1A",x"1A",x"C4",x"D5",x"B2",x"66",x"00",x"26",x"91",x"45",x"19",x"50",x"58",x"41",x"2B",x"80",x"D4",x"E3",x"BF",x"59",x"35",x"41",x"49",x"C8",x"C9",x"0B",x"CC",x"B0",x"6B",x"17",x"1A",x"3F",x"18",x"5B",x"E8",x"43",x"A0",x"9C",x"08",x"2F",x"4C",x"4B",x"47",x"95",x"36",x"E4",x"DC",x"44",x"33",x"CC",x"C2",x"48",x"01",x"86",x"17",x"D2",x"32",x"DD",x"04",x"C9",x"C8",x"05",x"24",x"75",x"C5",x"11",x"AA",x"25",x"A3",x"5B",x"76",x"CD",x"DA",x"AB",x"63",x"76",x"11",x"DB",x"92",x"04",x"6F",x"64",x"A7",x"CC",x"6A",x"5E",x"ED",x"47",x"EA",x"8D",x"B8",x"0B",x"30",x"2A",x"79",x"02",x"DF",x"CF",x"A5",x"02",x"A6",x"03",x"FD",x"28",x"03",x"A5",x"F2",x"6B",x"3A",x"BA",x"2A",x"22",x"95",x"92",x"BF",x"94",x"61",x"4F",x"08",x"51",x"BE",x"29",x"4A",x"15",x"04",x"28",x"D8",x"4A",x"D8",x"06",x"0E",x"4E",x"05",x"01",x"2D",x"46",x"38",x"E9",x"50",x"ED",x"85",x"2E",x"29",x"22",x"9F",x"39",x"91",x"64",x"68",x"22",x"AA",x"A0",x"2C",x"A3",x"97",x"CD",x"61",x"07",x"65",x"73",x"A2",x"48",x"B4",x"A5",x"12",x"05",x"8E",x"6F",x"17",x"0C",x"4C",x"22",x"11",x"2B",x"19",x"05",x"8B",x"2B",x"2E",x"5E",x"20",x"D4",x"77",x"6A",x"2F",x"10",x"74",x"51",x"5F",x"D0",x"62",x"54",x"B8",x"A6",x"7D",x"1A",x"1A",x"96",x"28",x"54",x"58",x"EC",x"1B",x"E1",x"89",x"02",x"8A",x"1F",x"14",x"A2",x"1C",x"3C",x"15",x"B8",x"57",x"20",x"5B",x"47",x"1C",x"42",x"93",x"02",x"0F",x"1D",x"57",x"0A",x"8A",x"A4",x"05",x"C0",x"80",x"FC",x"1E",x"87",x"28",x"06",x"55",x"50",x"70",x"8E",x"62",x"1F",x"90",x"02",x"E8",x"18",x"9F",x"AF",x"CA",x"14",x"CB",x"05",x"11",x"74",x"D3",x"ED",x"71",x"20",x"B8",x"4A",x"38",x"AE",x"1E",x"63",x"41",x"34",x"90",x"62",x"71",x"81",x"CF",x"39",x"C4",x"70",x"87",x"F5",x"32",x"5B",x"2E",x"32",x"02",x"CB",x"26",x"FD",x"A2",x"0C",x"AD",x"9F",x"4B",x"77",x"CB",x"37",x"39",x"17",x"2D",x"E7",x"5D",x"8A",x"2B",x"98",x"0D",x"6F",x"6F",x"33",x"73",x"AA",x"F0",x"0A",x"65",x"BF",x"8A",x"4C",x"C5",x"B0",x"4A",x"9B",x"06",x"E2",x"A9",x"88",x"31",x"32",x"E2",x"49",x"05",x"7A",x"F1",x"12",x"08",x"15",x"0E",x"15",x"04",x"09",x"A9",x"CB",x"88",x"9E",x"14",x"25",x"92",x"09",x"4F",x"B1",x"CB",x"08",x"63",x"92",x"B2",x"AE",x"29",x"6E",x"24",x"29",x"57",x"87",x"72",x"36",x"67",x"4C",x"51",x"BC",x"7B",x"A8",x"4A",x"44",x"49",x"8C",x"3C",x"D0",x"38",x"7F",x"C7",x"05",x"8A",x"9B",x"77",x"8C",x"32",x"D5",x"E8",x"CF",x"9C",x"78",x"65",x"50",x"E0",x"85",x"85",x"11",x"91",x"BA",x"3C",x"89",x"10",x"8F",x"90",x"88",x"0B",x"C3",x"57",x"6A",x"01",x"1E",x"36",x"0A",x"C8",x"52",x"E3",x"30",x"4A",x"53",x"D4",x"08",x"75",x"90",x"09",x"BB",x"49",x"4C",x"7F",x"52",x"E5",x"17",x"B1",x"D6",x"D9",x"F3",x"8A",x"09",x"99",x"62",x"E9",x"69",x"69",x"89",x"6D",x"3D",x"38",x"9F",x"81",x"06",x"8A",x"97",x"34",x"09",x"7C",x"09",x"60",x"05",x"09",x"BC",x"09",x"80",x"ED",x"94",x"80",x"9F",x"EB",x"01",x"FB",x"0E",x"3A",x"00",x"38",x"10",x"F8",x"68",x"03",x"4A",x"C3",x"4E",x"4C",x"7F",x"4F",x"B6",x"9A",x"0C",x"C8",x"B7",x"13",x"01",x"50",x"64",x"66",x"17",x"00",x"DA",x"72",x"00",x"03",x"6F",x"AD",x"03",x"62",x"3B",x"78",x"6E",x"2A",x"D6",x"80",x"6A",x"E7",x"EF",x"95",x"61",x"C9",x"01",x"F5",x"12",x"26",x"6D",x"5D",x"EA",x"6B",x"A2",x"A1",x"C1",x"07",x"53",x"B5",x"12",x"20",x"13",x"D0",x"53",x"DD",x"6B",x"A0",x"0D",x"C1",x"4E",x"2D",x"2F",x"1B",x"A0",x"03",x"A1",x"57",x"07",x"AD",x"3D",x"78",x"9E",x"44",x"DA",x"71",x"C0",x"AC",x"33",x"8A",x"67",x"B8",x"40",x"2A",x"BA",x"4E",x"4F",x"86",x"AE",x"2A",x"95",x"3F",x"64",x"EB",x"2D",x"79",x"D6",x"6C",x"23",x"3A",x"E8",x"03",x"F4",x"C0",x"03",x"19",x"A7",x"B0",x"7D",x"E4",x"DE",x"02",x"C4",x"2B",x"A5",x"F1",x"72",x"C9",x"00",x"8A",x"E9",x"7C",x"50",x"28",x"49",x"80",x"10",x"EB",x"38",x"C8",x"37",x"79",x"2C",x"AF",x"4B",x"2B",x"9C",x"CA",x"53",x"D0",x"67",x"61",x"CB",x"93",x"7D",x"85",x"F7",x"61",x"A7",x"0A",x"CE",x"AB",x"38",x"0B",x"F9",x"EA",x"3C",x"DC",x"20",x"97",x"61",x"80",x"F3",x"B5",x"A0",x"57",x"8E",x"84",x"C2",x"12",x"27",x"F0",x"7B",x"EA",x"AE",x"75",x"F5",x"00",x"64",x"84",x"01",x"18",x"23",x"15",x"70",x"D0",x"42",x"60",x"75",x"FE",x"8D",x"4B",x"28",x"6B",x"76",x"B5",x"CD",x"04",x"2B",x"A8",x"53",x"10",x"0E",x"D1",x"80",x"1C",x"E7",x"2F",x"71",x"0E",x"27",x"45",x"39",x"02",x"35",x"08",x"A9",x"53",x"92",x"5C",x"09",x"47",x"54",x"82",x"D3",x"A2",x"09",x"32",x"6B",x"36",x"01",x"21",x"88",x"BA",x"A4",x"44",x"5F",x"93",x"9C",x"2D",x"95",x"B6",x"AA",x"62",x"AD",x"0F",x"5A",x"88",x"58",x"95",x"03",x"5B",x"68",x"0B",x"F8",x"0B",x"C0",x"0A",x"0B",x"02",x"88",x"0B",x"70",x"02",x"A1",x"51",x"51",x"2A",x"D0",x"61",x"AA",x"7F",x"68",x"4C",x"70",x"C4",x"95",x"50",x"5B",x"D1",x"80",x"B5",x"32",x"EB",x"29",x"0F",x"57",x"23",x"21",x"4D",x"B8",x"B8",x"0F",x"C6",x"12",x"03",x"04",x"80",x"2A",x"1F",x"AF",x"4F",x"21",x"0B",x"1E",x"35",x"63",x"65",x"F0",x"0E",x"5F",x"61",x"06",x"80",x"0C",x"78",x"57",x"B7",x"86",x"B7",x"B4",x"AE",x"40",x"E7",x"0A",x"D0",x"F0",x"04",x"46",x"04",x"01",x"09",x"A2",x"71",x"98",x"E6",x"09",x"99",x"34",x"33",x"E2",x"E5",x"96",x"F6",x"FA",x"76",x"20",x"6C",x"64",x"9C",x"D8",x"4F",x"BA",x"0C",x"CE",x"4F",x"91",x"7C",x"00",x"AE",x"60",x"17",x"81",x"CE",x"4C",x"BC",x"D3",x"EF",x"85",x"62",x"3D",x"29",x"39",x"37",x"07",x"F1",x"9E",x"E0",x"2F",x"38",x"17",x"89",x"9C",x"B1",x"C2",x"A0",x"AA",x"31",x"55",x"47",x"E3",x"F5",x"29",x"BB",x"90",x"B7",x"FB",x"04",x"52",x"AC",x"EE",x"2C",x"70",x"AA",x"4C",x"12",x"F8",x"A8",x"98",x"3C",x"00",x"52",x"A6",x"A4",x"81",x"0E",x"A4",x"22",x"A7",x"26",x"22",x"85",x"91",x"08",x"22",x"2F",x"87",x"EA",x"5D",x"90",x"FF",x"B1",x"0F",x"AE",x"35",x"5D",x"38",x"07",x"79",x"15",x"DC",x"27",x"15",x"00",x"4E",x"42",x"EE",x"1C",x"9A",x"CC",x"21",x"65",x"B1",x"61",x"8D",x"40",x"80",x"AF",x"1C",x"39",x"10",x"D1",x"13",x"2F",x"F0",x"01",x"8C",x"C8",x"20",x"6E",x"64",x"7F",x"3A",x"A0",x"44",x"92",x"4A",x"DE",x"18",x"D4",x"DC",x"D9",x"F4",x"4C",x"9F",x"6A",x"4C",x"2B",x"A5",x"EE",x"B0",x"E0",x"AE",x"CA",x"51",x"A2",x"96",x"7B",x"98",x"A9",x"C2",x"10",x"80",x"3E",x"EB",x"0A",x"25",x"DE",x"05",x"68",x"CC",x"A2",x"C6",x"7E",x"C8",x"A2",x"75",x"4F",x"21",x"A9",x"6F",x"71",x"C4",x"87",x"50",x"C0",x"32",x"4A",x"35",x"17",x"6D",x"03",x"EC",x"9E",x"0B",x"47",x"42",x"9C",x"6A",x"07",x"30",x"02",x"29",x"C3",x"01",x"69",x"DD",x"C0",x"A4",x"A2",x"58",x"6B",x"AD",x"8F",x"F0",x"FB",x"8D",x"FD",x"9C",x"10",x"D8",x"D6",x"05",x"DD",x"2C",x"79",x"60",x"F4",x"40",x"86",x"09",x"00",x"36",x"6B",x"01",x"D8",x"94",x"86",x"85",x"3C",x"D6",x"A0",x"8D",x"2C",x"8E",x"B7",x"A2",x"04",x"2F",x"A5",x"35",x"59",x"8C",x"2D",x"D4",x"80",x"2E",x"4B",x"4E",x"C2",x"A1",x"84",x"8F",x"B4",x"AF",x"A9",x"A9",x"CA",x"95",x"67",x"A4",x"56",x"6A",x"66",x"A3",x"24",x"35",x"33",x"79",x"49",x"AD",x"A1",x"7D",x"BF",x"9C",x"05",x"19",x"97",x"60",x"6C",x"89",x"0C",x"C2",x"7A",x"8E",x"41",x"61",x"D4",x"AC",x"5B",x"8F",x"8F",x"80",x"1D",x"5C",x"90",x"1D",x"AD",x"12",x"D0",x"D2",x"02",x"F9",x"F0",x"F9",x"83",x"D7",x"1C",x"8E",x"81",x"17",x"23",x"36",x"67",x"4B",x"DF",x"63",x"D7",x"DC",x"41",x"75",x"99",x"D1",x"52",x"C3",x"B7",x"08",x"9C",x"64",x"3B",x"A0",x"01",x"5E",x"B9",x"34",x"86",x"B7",x"29",x"35",x"AB",x"2D",x"90",x"41",x"DA",x"39",x"A4",x"FF",x"49",x"B8",x"C5",x"8A",x"AC",x"95",x"64",x"34",x"5B",x"67",x"F0",x"EB",x"1C",x"0D",x"11",x"8A",x"A6",x"4F",x"36",x"6F",x"6D",x"41",x"21",x"53",x"6A",x"42",x"01",x"4B",x"57",x"90",x"D2",x"A8",x"42",x"14",x"D1",x"92",x"42",x"14",x"D0",x"92",x"AD",x"CF",x"D2",x"78",x"5B",x"CD",x"6F",x"65",x"AE",x"4A",x"94",x"92",x"B1",x"0B",x"43",x"31",x"EA",x"10",x"C5",x"27",x"1B",x"62",x"A8",x"16",x"E8",x"03",x"DE",x"06",x"86",x"21",x"53",x"07",x"39",x"C9",x"64",x"C9",x"8A",x"04",x"CB",x"61",x"AB",x"E9",x"00",x"B0",x"EE",x"CD",x"05",x"A0",x"08",x"7E",x"F7",x"28",x"20",x"B3",x"C9",x"64",x"05",x"D3",x"53",x"64",x"80",x"B1",x"04",x"A9",x"40",x"A2",x"76",x"A8",x"5F",x"3D",x"5F",x"E0",x"D2",x"C3",x"32",x"BA",x"0D",x"B6",x"AE",x"B1",x"2B",x"E7",x"BF",x"0A",x"4D",x"82",x"AF",x"60",x"2C",x"85",x"F4",x"4E",x"89",x"69",x"36",x"9D",x"21",x"65",x"D6",x"2C",x"4B",x"9A",x"05",x"6B",x"92",x"81",x"A6",x"21",x"1B",x"1A",x"D0",x"C7",x"1D",x"08",x"8A",x"17",x"02",x"36",x"04",x"34",x"AD",x"99",x"6D",x"AE",x"9A",x"75",x"E9",x"18",x"69",x"E8",x"AB",x"9C",x"47",x"9C",x"1F",x"65",x"A5",x"05",x"F8",x"9E",x"4C",x"BC",x"55",x"7B",x"3F",x"43",x"A9",x"28",x"F0",x"80",x"1A",x"07",x"37",x"C7",x"A8",x"00",x"4D",x"B1",x"CB",x"53",x"09",x"A8",x"BB",x"92",x"0A",x"A2",x"EE",x"C3",x"A9",x"50",x"AF",x"20",x"8E",x"9F",x"80",x"39",x"5D",x"21",x"38",x"E9",x"01",x"8D",x"7F",x"CC",x"54",x"CE",x"5B",x"AD",x"A5",x"6C",x"0D",x"A6",x"7D",x"E9",x"D0",x"37",x"C7",x"55",x"DD",x"27",x"04",x"40",x"D0",x"7C",x"BF",x"38",x"C9",x"01",x"F0",x"6C",x"FC",x"05",x"03",x"D0",x"C1",x"B7",x"98",x"2B",x"61",x"0B",x"97",x"6B",x"B3",x"B2",x"0A",x"29",x"E8",x"67",x"D0",x"2C",x"20",x"F0",x"62",x"7F",x"96",x"25",x"05",x"6C",x"95",x"85",x"AD",x"AE",x"AD",x"94",x"AD",x"A5",x"93",x"75",x"D7",x"20",x"9D",x"6A",x"A9",x"F6",x"AF",x"9D",x"79",x"46",x"04",x"64",x"05",x"67",x"9B",x"6A",x"A2",x"85",x"5D",x"5C",x"9F",x"A6",x"2C",x"80",x"87",x"AD",x"16",x"1A",x"29",x"0F",x"8D",x"FB",x"D0",x"20",x"B5",x"E8",x"4A",x"91",x"18",x"A9",x"01",x"47",x"1D",x"3D",x"A0",x"04",x"B1",x"02",x"F2",x"0F",x"03",x"93",x"AB",x"54",x"D4",x"1F",x"6A",x"CE",x"55",x"62",x"80",x"71",x"AC",x"AA",x"46",x"82",x"F5",x"58",x"25",x"19",x"BA",x"2F",x"F6",x"0A",x"CE",x"E4",x"60",x"3C",x"7C",x"B6",x"B4",x"BB",x"EE",x"CC",x"4E",x"47",x"45",x"48",x"CA",x"E4",x"2D",x"29",x"6B",x"52",x"46",x"08",x"6C",x"D6",x"D7",x"A0",x"D5",x"01",x"84",x"9E",x"AD",x"03",x"28",x"88",x"14",x"92",x"08",x"34",x"F0",x"A0",x"E0",x"FF",x"3F",x"25",x"02",x"18",x"30",x"22",x"28",x"53",x"20",x"E0",x"E8",x"C3",x"38",x"46",x"78",x"48",x"58",x"D8",x"C0",x"FF",x"6F",x"53",x"66",x"24",x"5A",x"74",x"93",x"AB",x"A6",x"A8",x"F8",x"E0",x"F5",x"81",x"57",x"4D",x"FC",x"7C",x"D1",x"1C",x"04",x"1F",x"6E",x"8A",x"A8",x"A4",x"70",x"0D",x"07",x"98",x"C0",x"6C",x"77",x"56",x"1C",x"22",x"C2",x"58",x"44",x"34",x"88",x"70",x"9F",x"20",x"3A",x"02",x"FD",x"4C",x"54",x"54",x"E9",x"F6",x"3A",x"79",x"35",x"2A",x"52",x"36",x"4F",x"28",x"94",x"74",x"0C",x"08",x"58",x"EC",x"3A",x"CA",x"60",x"20",x"86",x"CE",x"57",x"5C",x"08",x"75",x"9B",x"CD",x"28",x"6F",x"A6",x"24",x"2B",x"06",x"45",x"4D",x"FE",x"7C",x"2B",x"57",x"64",x"87",x"AA",x"02",x"B0",x"AB",x"CB",x"0D",x"16",x"80",x"24",x"40",x"FE",x"42",x"76",x"2B",x"7C",x"FD",x"1E",x"F8",x"79",x"C4",x"0F",x"E9",x"8C",x"8C",x"5E",x"78",x"92",x"70",x"CE",x"CC",x"7E",x"5F",x"06",x"FF",x"A6",x"42",x"4C",x"08",x"64",x"B0",x"A9",x"26",x"B7",x"C9",x"C7",x"4C",x"FE",x"A1",x"04",x"48",x"E8",x"C8",x"31",x"0C",x"60",x"47",x"B3",x"0A",x"80",x"31",x"94",x"04",x"F9",x"BB",x"C0",x"80",x"F9",x"AC",x"FC",x"EC",x"F9",x"2C",x"70",x"13",x"67",x"0E",x"38",x"60",x"C4",x"7F",x"C9",x"51",x"73",x"33",x"1C",x"3C",x"D4",x"CC",x"FE",x"17",x"7B",x"86",x"0C",x"0C",x"8C",x"FA",x"63",x"A5",x"EA",x"BC",x"7F",x"92",x"78",x"DA",x"08",x"E6",x"AB",x"A9",x"DA",x"50",x"6E",x"36",x"87",x"E2",x"63",x"52",x"84",x"98",x"31",x"AC",x"09",x"33",x"C3",x"04",x"8B",x"DC",x"30",x"8B",x"0C",x"73",x"10",x"9F",x"49",x"67",x"32",x"34",x"4E",x"53",x"76",x"0F",x"F8",x"67",x"D1",x"B8",x"A2",x"1A",x"CE",x"8E",x"1C",x"8C",x"E8",x"34",x"67",x"08",x"8B",x"2A",x"78",x"67",x"11",x"11",x"3C",x"F8",x"D7",x"8C",x"70",x"9E",x"36",x"01",x"BB",x"5B",x"C0",x"63",x"04",x"F8",x"67",x"88",x"07",x"D5",x"EC",x"7C",x"2E",x"04",x"AF",x"0A",x"8E",x"CF",x"3D",x"67",x"C3",x"02",x"63",x"1F",x"43",x"31",x"0D",x"CC",x"5C",x"0C",x"2C",x"E0",x"67",x"B1",x"50",x"80",x"4B",x"64",x"0C",x"67",x"14",x"0D",x"35",x"ED",x"04",x"FF",x"C0",x"60",x"30",x"62",x"8F",x"5F",x"06",x"2D",x"6E",x"8A",x"B7",x"85",x"84",x"16",x"50",x"8E",x"78",x"0C",x"97",x"30",x"EA",x"0E",x"18",x"B1",x"26",x"36",x"97",x"8C",x"E9",x"43",x"6C",x"E6",x"93",x"74",x"CC",x"87",x"F4",x"0D",x"18",x"DE",x"9C",x"D1",x"16",x"78",x"6C",x"FD",x"41",x"38",x"BA",x"6F",x"3E",x"C6",x"7F",x"6B",x"35",x"63",x"E8",x"45",x"51",x"0C",x"9F",x"18",x"25",x"48",x"87",x"7C",x"B5",x"18",x"09",x"45",x"06",x"2A",x"60",x"44",x"05",x"65",x"18",x"3E",x"9A",x"EF",x"6F",x"06",x"F7",x"53",x"42",x"7E",x"09",x"0E",x"91",x"87",x"31",x"99",x"8F",x"A2",x"D9",x"41",x"63",x"6B",x"7F",x"3E",x"36",x"FE",x"61",x"18",x"A2",x"3C",x"A7",x"19",x"87",x"A1",x"46",x"35",x"51",x"0D",x"AF",x"DE",x"4F",x"63",x"28",x"64",x"40",x"B0",x"4D",x"5A",x"95",x"60",x"0C",x"D7",x"0D",x"1E",x"32",x"92",x"F6",x"EB",x"2B",x"45",x"0A",x"82",x"B0",x"FE",x"0F",x"02",x"DC",x"FA",x"21",x"CF",x"7E",x"0C",x"81",x"50",x"35",x"47",x"0D",x"D4",x"4E",x"44",x"AB",x"B9",x"99",x"03",x"31",x"9D",x"CC",x"AF",x"BB",x"34",x"D5",x"AD",x"03",x"44",x"7C",x"3E",x"35",x"CC",x"9C",x"7D",x"32",x"A2",x"B3",x"04",x"0C",x"94",x"90",x"7C",x"48",x"F0",x"D8",x"F4",x"87",x"00",x"C0",x"4C",x"AA",x"3D",x"EE",x"5A",x"90",x"D6",x"16",x"BA",x"34",x"32",x"DC",x"ED",x"B0",x"0B",x"B7",x"02",x"D8",x"07",x"D7",x"0B",x"14",x"09",x"D4",x"D8",x"6C",x"57",x"39",x"F8",x"9A",x"1B",x"A2",x"ED",x"C0",x"E0",x"78",x"0E",x"1C",x"F8",x"7D",x"1B",x"60",x"9E",x"1D",x"86",x"64",x"9E",x"58",x"5D",x"0F",x"91",x"49",x"D6",x"12",x"FE",x"EE",x"C6",x"FA",x"41",x"90",x"B1",x"84",x"81",x"A1",x"DC",x"78",x"7C",x"68",x"88",x"18",x"BC",x"30",x"EC",x"EB",x"85",x"00",x"86",x"15",x"FD",x"10",x"2A",x"80",x"18",x"47",x"89",x"12",x"7C",x"0A",x"90",x"9B",x"4D",x"FE",x"7E",x"20",x"74",x"40",x"C1",x"6A",x"03",x"AC",x"2B",x"3A",x"44",x"48",x"39",x"D9",x"40",x"F6",x"70",x"F0",x"26",x"60",x"FC",x"74",x"31",x"09",x"24",x"5A",x"7A",x"44",x"82",x"44",x"6C",x"DE",x"72",x"03",x"E3",x"72",x"18",x"64",x"90",x"73",x"2C",x"98",x"5B",x"72",x"5D",x"CD",x"8B",x"A2",x"B2",x"F1",x"8B",x"C0",x"08",x"D9",x"A8",x"38",x"A9",x"C5",x"4C",x"51",x"59",x"62",x"30",x"7C",x"04",x"2B",x"60",x"2A",x"8A",x"6A",x"82",x"B2",x"AA",x"44",x"2E",x"20",x"38",x"01",x"73",x"A9",x"20",x"6C",x"82",x"95",x"70",x"40",x"CA",x"C3",x"04",x"A4",x"B6",x"82",x"08",x"09",x"72",x"24",x"38",x"24",x"DB",x"CA",x"7C",x"42",x"E8",x"68",x"03",x"28",x"F6",x"40",x"00",x"0A",x"C2",x"18",x"04",x"7D",x"35",x"09",x"60",x"E2",x"1D",x"9F",x"62",x"12",x"C4",x"30",x"14",x"30",x"85",x"8B",x"12",x"24",x"9E",x"0E",x"53",x"26",x"2F",x"42",x"C4",x"48",x"E4",x"56",x"22",x"8F",x"86",x"B6",x"C2",x"44",x"C8",x"52",x"E6",x"4A",x"84",x"FE",x"C1",x"6A",x"60",x"B6",x"90",x"1C",x"92",x"43",x"71",x"ED",x"0E",x"05",x"D0",x"3B",x"14",x"64",x"98",x"5F",x"28",x"48",x"42",x"10",x"C7",x"40",x"30",x"29",x"FC",x"CC",x"E4",x"3E",x"A6",x"28",x"4E",x"D0",x"88",x"8E",x"D3",x"AD",x"A9",x"C0",x"86",x"3A",x"40",x"D1",x"AB",x"1D",x"8C",x"AB",x"1D",x"8A",x"AB",x"1D",x"0A",x"A8",x"05",x"60",x"7C",x"E4",x"DB",x"0E",x"C6",x"6D",x"87",x"42",x"32",x"14",x"69",x"2B",x"AE",x"12",x"AC",x"EC",x"C8",x"42",x"F8",x"7B",x"22",x"94",x"68",x"58",x"48",x"F4",x"BB",x"1D",x"8C",x"C7",x"1D",x"8A",x"A9",x"1D",x"28",x"8A",x"50",x"0F",x"45",x"B3",x"09",x"58",x"DD",x"BE",x"92",x"29",x"9A",x"44",x"B2",x"3F",x"1A",x"AD",x"2C",x"34",x"24",x"58",x"F4",x"3F",x"72",x"60",x"20",x"BC",x"28",x"CE",x"56",x"1C",x"1A",x"60",x"8D",x"78",x"3D",x"DA",x"6C",x"38",x"FC",x"95",x"90",x"F8",x"42",x"CC",x"FC",x"83",x"C0",x"C6",x"26",x"10",x"64",x"68",x"68",x"A4",x"A4",x"20",x"71",x"10",x"F1",x"60",x"FC",x"5C",x"0C",x"3D",x"48",x"0F",x"46",x"DE",x"78",x"08",x"8E",x"CC",x"7C",x"7E",x"24",x"EC",x"32",x"87",x"90",x"9E",x"BA",x"09",x"58",x"32",x"20",x"D1",x"4B",x"72",x"28",x"B0",x"76",x"51",x"60",x"7C",x"D9",x"03",x"F1",x"69",x"7E",x"60",x"3C",x"7E",x"20",x"0F",x"86",x"6D",x"87",x"42",x"3A",x"14",x"7E",x"73",x"06",x"4C",x"6A",x"20",x"50",x"D1",x"12",x"24",x"18",x"F4",x"89",x"7C",x"E9",x"22",x"CF",x"58",x"87",x"E2",x"B6",x"10",x"C5",x"83",x"14",x"28",x"B1",x"61",x"A6",x"47",x"32",x"F9",x"3C",x"90",x"C0",x"06",x"7C",x"64",x"D4",x"80",x"55",x"3A",x"4C",x"54",x"64",x"B8",x"FF",x"6A",x"07",x"20",x"46",x"D6",x"A1",x"10",x"28",x"F8",x"A0",x"44",x"58",x"01",x"C6",x"7E",x"64",x"08",x"10",x"D7",x"17",x"05",x"8B",x"92",x"48",x"A0",x"70",x"40",x"87",x"24",x"6C",x"96",x"3E",x"0C",x"CF",x"78",x"35",x"C4",x"20",x"17",x"62",x"B3",x"AA",x"96",x"F0",x"E3",x"5C",x"69",x"DE",x"D0",x"55",x"8E",x"7C",x"AA",x"60",x"57",x"6E",x"A6",x"D0",x"6A",x"3A",x"C9",x"B3",x"B2",x"8D",x"A2",x"95",x"B1",x"5F",x"A9",x"6D",x"A2",x"CD",x"D8",x"20",x"80",x"FC",x"31",x"A5",x"93",x"3A",x"16",x"FE",x"67",x"17",x"60",x"F9",x"11",x"94",x"43",x"98",x"62",x"AD",x"54",x"FB",x"DA",x"15",x"1E",x"3D",x"62",x"CE",x"0F",x"28",x"EC",x"75",x"20",x"09",x"5E",x"72",x"5E",x"65",x"18",x"B2",x"16",x"B8",x"A4",x"0A",x"9D",x"84",x"0B",x"8F",x"38",x"BB",x"E9",x"30",x"90",x"2C",x"C9",x"BF",x"B0",x"28",x"35",x"E6",x"48",x"C8",x"95",x"19",x"0C",x"C5",x"54",x"48",x"CC",x"2C",x"AE",x"CC",x"29",x"68",x"9E",x"65",x"23",x"58",x"90",x"D1",x"E6",x"F7",x"B0",x"CD",x"ED",x"EA",x"8B",x"AC",x"28",x"61",x"A1",x"99",x"39",x"51",x"60",x"A9",x"BB",x"EF",x"7B",x"18",x"6D",x"CB",x"F4",x"3D",x"2A",x"06",x"29",x"76",x"A6",x"1B",x"4C",x"8F",x"20",x"F3",x"DA",x"5D",x"B4",x"2B",x"F8",x"B1",x"EE",x"97",x"BC",x"F3",x"A7",x"66",x"94",x"5E",x"DE",x"D8",x"68",x"13",x"50",x"AE",x"B9",x"CF",x"0A",x"3E",x"4A",x"4C",x"CE",x"3A",x"0A",x"82",x"67",x"C3",x"84",x"5B",x"18",x"66",x"20",x"DE",x"86",x"5E",x"EC",x"5B",x"C3",x"67",x"48",x"B9",x"4D",x"B9",x"FB",x"00",x"99",x"7A",x"D3",x"88",x"10",x"F7",x"68",x"7D",x"16",x"17",x"AD",x"18",x"27",x"19",x"E0",x"53",x"78",x"58",x"86",x"1B",x"59",x"AB",x"A5",x"91",x"94",x"50",x"CE",x"8A",x"7E",x"8D",x"51",x"79",x"F2",x"E9",x"A5",x"F4",x"B6",x"85",x"2C",x"F8",x"18",x"CC",x"0B",x"D1",x"94",x"2D",x"43",x"F5",x"9B",x"CB",x"D0",x"F1",x"98",x"5E",x"65",x"A3",x"18",x"E8",x"8A",x"C2",x"38",x"B4",x"0A",x"56",x"A5",x"AD",x"19",x"E5",x"0B",x"85",x"0D",x"BF",x"0C",x"F0",x"25",x"20",x"F5",x"D6",x"62",x"A0",x"05",x"5F",x"1B",x"1A",x"CF",x"0B",x"F3",x"0A",x"24",x"0D",x"98",x"52",x"D7",x"0C",x"89",x"F4",x"89",x"4F",x"48",x"FE",x"E8",x"5D",x"AA",x"7E",x"EC",x"A2",x"05",x"BD",x"A8",x"7F",x"95",x"16",x"FE",x"55",x"F8",x"60",x"BB",x"30",x"20",x"25",x"E4",x"A5",x"F6",x"5D",x"E2",x"BD",x"79",x"89",x"2C",x"0B",x"9D",x"2F",x"CA",x"10",x"FA",x"3B",x"27",x"2D",x"B2",x"AF",x"19",x"BC",x"2B",x"B5",x"B0",x"10",x"BC",x"20",x"B5",x"05",x"BA",x"2A",x"46",x"07",x"23",x"D6",x"A9",x"15",x"4E",x"B0",x"93",x"9A",x"5F",x"61",x"C9",x"30",x"DD",x"F2",x"28",x"31",x"8E",x"B3",x"C4",x"7F",x"5D",x"0C",x"DC",x"5F",x"B4",x"9F",x"5E",x"B5",x"56",x"D8",x"8C",x"45",x"41",x"2E",x"1B",x"AC",x"10",x"F2",x"41",x"2A",x"D6",x"78",x"38",x"F2",x"88",x"4C",x"FE",x"F4",x"3E",x"D5",x"C0",x"8E",x"5D",x"5F",x"B1",x"18",x"77",x"5A",x"19",x"AD",x"48",x"B5",x"15",x"54",x"D6",x"11",x"5A",x"4A",x"47",x"08",x"CC",x"EB",x"0E",x"4C",x"99",x"ED",x"93",x"D0",x"B8",x"A4",x"C6",x"4C",x"09",x"2C",x"FC",x"BA",x"F6",x"BB",x"92",x"CF",x"86",x"26",x"B1",x"61",x"EC",x"5D",x"5D",x"43",x"33",x"9D",x"C0",x"06",x"6E",x"B2",x"F0",x"35",x"D4",x"44",x"0B",x"31",x"49",x"D0",x"2D",x"79",x"00",x"B1",x"AD",x"86",x"20",x"AD",x"B0",x"39",x"68",x"02",x"A2",x"2B",x"8E",x"9F",x"CC",x"47",x"A4",x"05",x"30",x"0B",x"AC",x"B9",x"FE",x"45",x"8C",x"BB",x"B2",x"EE",x"BA",x"7F",x"F4",x"0A",x"BA",x"88",x"4E",x"B1",x"15",x"72",x"88",x"92",x"6A",x"10",x"C8",x"B1",x"1A",x"E4",x"56",x"3F",x"BB",x"C9",x"4F",x"E4",x"BB",x"41",x"20",x"5E",x"AC",x"27",x"4A",x"17",x"48",x"19",x"BE",x"87",x"04",x"97",x"06",x"E2",x"24",x"68",x"C4",x"08",x"5A",x"C1",x"6F",x"50",x"88",x"D0",x"EA",x"65",x"B8",x"A9",x"E8",x"8E",x"D3",x"36",x"A9",x"3B",x"27",x"B8",x"C9",x"53",x"BB",x"0C",x"20",x"32",x"5E",x"8D",x"FE",x"8E",x"E5",x"9B",x"C5",x"55",x"D0",x"0B",x"FC",x"0A",x"54",x"11",x"1C",x"C1",x"26",x"DA",x"C9",x"D8",x"D0",x"EF",x"29",x"48",x"AD",x"B2",x"CF",x"67",x"0A",x"30",x"2B",x"41",x"A9",x"D8",x"7C",x"AE",x"52",x"15",x"25",x"A0",x"84",x"F5",x"CE",x"5E",x"68",x"C9",x"58",x"7A",x"7D",x"9F",x"85",x"31",x"6B",x"2A",x"2C",x"61",x"7D",x"94",x"AD",x"CF",x"2C",x"AE",x"D0",x"5D",x"20",x"4B",x"6B",x"8D",x"3D",x"68",x"8E",x"D2",x"37",x"3B",x"0D",x"AC",x"F0",x"B2",x"15",x"AE",x"B6",x"17",x"EC",x"5D",x"AD",x"B7",x"F6",x"A8",x"68",x"C7",x"06",x"8E",x"9C",x"8C",x"D8",x"C6",x"38",x"B4",x"56",x"C3",x"D1",x"4E",x"AA",x"AD",x"33",x"ED",x"D2",x"FB",x"EC",x"95",x"C2",x"E3",x"B5",x"95",x"FF",x"15",x"8D",x"95",x"B4",x"A5",x"D0",x"52",x"62",x"A9",x"6A",x"AD",x"AF",x"7F",x"EB",x"BF",x"20",x"BE",x"9E",x"5E",x"4C",x"0E",x"5F",x"BF",x"D3",x"52",x"42",x"B3",x"D4",x"7F",x"3E",x"9C",x"07",x"CD",x"F9",x"7C",x"18",x"98",x"65",x"17",x"DB",x"77",x"20",x"68",x"A9",x"AC",x"E2",x"00",x"C6",x"21",x"30",x"0E",x"32",x"71",x"D0",x"38",x"08",x"39",x"0C",x"05",x"15",x"9E",x"06",x"CC",x"0A",x"18",x"B9",x"1A",x"EC",x"9E",x"C0",x"DA",x"85",x"A6",x"DB",x"AA",x"6F",x"A0",x"45",x"F4",x"8F",x"06",x"75",x"FF",x"E0",x"80",x"B0",x"02",x"3E",x"3E",x"16",x"38",x"06",x"AA",x"D5",x"33",x"12",x"A0",x"76",x"52",x"EA",x"53",x"85",x"AD",x"98",x"54",x"AE",x"A5",x"55",x"79",x"77",x"6D",x"CC",x"AB",x"25",x"DE",x"F7",x"AE",x"67",x"77",x"AC",x"A7",x"E3",x"E3",x"35",x"15",x"92",x"C5",x"8D",x"76",x"90",x"EC",x"05",x"01",x"4A",x"18",x"29",x"0F",x"F2",x"BD",x"AF",x"82",x"76",x"3F",x"5F",x"38",x"F8",x"12",x"36",x"A4",x"15",x"27",x"5E",x"77",x"28",x"88",x"88",x"E2",x"C0",x"7A",x"04",x"F8",x"05",x"F0",x"06",x"E1",x"07",x"43",x"8A",x"17",x"E3",x"C3",x"CE",x"02",x"DB",x"AD",x"01",x"5D",x"B4",x"B1",x"18",x"BD",x"7B",x"79",x"F2",x"FC",x"E8",x"E0",x"08",x"EE",x"90",x"F6",x"60",x"8C",x"5F",x"98",x"2C",x"AD",x"49",x"2B",x"18",x"F3",x"0B",x"4B",x"68",x"90",x"AC",x"01",x"E8",x"0F",x"23",x"C1",x"89",x"4A",x"10",x"F9",x"F3",x"99",x"12",x"69",x"6C",x"AC",x"D5",x"5F",x"55",x"22",x"8D",x"8E",x"CF",x"86",x"0B",x"D4",x"38",x"01",x"D6",x"D2",x"A9",x"10",x"20",x"8C",x"61",x"AA",x"FD",x"47",x"C9",x"61",x"29",x"A1",x"F1",x"B6",x"FF",x"77",x"4A",x"AE",x"D1",x"24",x"A3",x"3B",x"E2",x"A2",x"09",x"0E",x"B7",x"9A",x"68",x"E0",x"0F",x"0E",x"C9",x"00",x"D0",x"7B",x"D6",x"0C",x"51",x"0A",x"C9",x"20",x"92",x"92",x"6C",x"1A",x"A3",x"18",x"C9",x"EC",x"B7",x"14",x"D6",x"AD",x"C4",x"5C",x"AD",x"D7",x"7F",x"40",x"FF",x"31",x"EE",x"09",x"ED",x"A6",x"D0",x"A5",x"4C",x"9F",x"69",x"FD",x"72",x"4C",x"65",x"20",x"DE",x"E4",x"6B",x"1F",x"C7",x"F2",x"E9",x"31",x"E8",x"C8",x"9C",x"8D",x"1C",x"8A",x"98",x"11",x"99",x"B4",x"0D",x"0B",x"E8",x"9D",x"D8",x"69",x"1A",x"2B",x"FD",x"05",x"37",x"1F",x"D0",x"64",x"C7",x"00",x"EE",x"18",x"05",x"90",x"F0",x"97",x"58",x"34",x"F5",x"A4",x"B9",x"C9",x"04",x"79",x"05",x"06",x"9E",x"07",x"27",x"41",x"49",x"AA",x"A7",x"61",x"CC",x"55",x"01",x"33",x"5B",x"11",x"95",x"25",x"A3",x"A6",x"D8",x"EA",x"2B",x"48",x"18",x"85",x"2D",x"49",x"38",x"8C",x"CA",x"40",x"8C",x"4A",x"11",x"2F",x"A5",x"18",x"31",x"63",x"1A",x"87",x"61",x"19",x"08",x"42",x"65",x"19",x"72",x"F0",x"37",x"1F",x"2B",x"82",x"5D",x"1E",x"55",x"89",x"6A",x"E6",x"8C",x"4D",x"10",x"AC",x"9C",x"6A",x"31",x"D4",x"2B",x"10",x"A9",x"86",x"88",x"1B",x"55",x"0E",x"B2",x"D0",x"03",x"18",x"87",x"8A",x"D9",x"A4",x"84",x"A7",x"B9",x"69",x"05",x"22",x"EB",x"04",x"59",x"0C",x"0D",x"0B",x"D0",x"73",x"A3",x"C5",x"0A",x"99",x"03",x"F0",x"F1",x"B0",x"03",x"B5",x"D4",x"92",x"0C",x"28",x"50",x"29",x"38",x"09",x"52",x"08",x"20",x"9A",x"64",x"28",x"DA",x"9A",x"4E",x"4C",x"61",x"5A",x"C2",x"E6",x"05",x"24",x"48",x"68",x"C3",x"88",x"AA",x"54",x"F6",x"A1",x"CD",x"B5",x"40",x"25",x"38",x"F4",x"7D",x"B0",x"0D",x"CA",x"E0",x"FF",x"BF",x"08",x"56",x"E4",x"A1",x"C6",x"25",x"DE",x"0C",x"1D",x"76",x"5D",x"12",x"45",x"35",x"95",x"05",x"2D",x"31",x"46",x"C2",x"AA",x"60",x"3D",x"91",x"2B",x"8F",x"A2",x"68",x"84",x"B9",x"14",x"E8",x"A9",x"7E",x"09",x"E8",x"63",x"FF",x"04",x"9D",x"2A",x"05",x"92",x"60",x"49",x"9A",x"68",x"E0",x"8C",x"70",x"66",x"C6",x"E0",x"38",x"58",x"56",x"46",x"14",x"9F",x"A4",x"15",x"DD",x"24",x"58",x"73",x"03",x"4C",x"66",x"B7",x"AF",x"73",x"77",x"06",x"D3",x"0E",x"2A",x"0E",x"0F",x"96",x"04",x"10",x"CE",x"13",x"48",x"E7",x"D3",x"87",x"84",x"6C",x"2D",x"AA",x"48",x"F9",x"46",x"15",x"0E",x"14",x"95",x"13",x"6A",x"8E",x"BA",x"36",x"0B",x"66",x"0A",x"90",x"17",x"18",x"3F",x"E4",x"85",x"0F",x"64",x"15",x"13",x"D5",x"10",x"5A",x"45",x"14",x"D5",x"56",x"65",x"1B",x"CE",x"A1",x"D4",x"6D",x"D5",x"75",x"11",x"18",x"11",x"AC",x"51",x"DA",x"B0",x"62",x"1B",x"EB",x"60",x"6F",x"03",x"64",x"05",x"49",x"90",x"BF",x"4D",x"FD",x"59",x"4C",x"01",x"64",x"58",x"BC",x"CA",x"C2",x"48",x"8A",x"20",x"BC",x"62",x"C2",x"FF",x"D9",x"46",x"C3",x"10",x"3A",x"C6",x"54",x"1E",x"85",x"06",x"86",x"07",x"3F",x"4D",x"08",x"BA",x"A4",x"75",x"9D",x"60",x"E8",x"09",x"A8",x"0E",x"08",x"E9",x"A6",x"B5",x"07",x"06",x"AB",x"60",x"F9",x"27",x"56",x"73",x"9C",x"CB",x"54",x"2E",x"0A",x"88",x"AD",x"2A",x"0B",x"B1",x"55",x"25",x"04",x"B6",x"AA",x"05",x"44",x"AB",x"9B",x"FD",x"10",x"21",x"18",x"DE",x"AA",x"0E",x"01",x"E4",x"B6",x"6B",x"55",x"07",x"42",x"EE",x"55",x"87",x"31",x"9E",x"54",x"5F",x"69",x"D6",x"E8",x"77",x"F9",x"29",x"1F",x"6E",x"18",x"20",x"E9",x"6A",x"76",x"F0",x"0E",x"AF",x"27",x"88",x"EA",x"C2",x"1C",x"C5",x"19",x"32",x"05",x"8B",x"A6",x"E8",x"64",x"7C",x"32",x"74",x"04",x"73",x"01",x"E6",x"D5",x"8B",x"BA",x"84",x"92",x"0B",x"61",x"64",x"6B",x"10",x"B2",x"F3",x"73",x"99",x"E8",x"AA",x"B0",x"10",x"33",x"21",x"73",x"99",x"A9",x"0A",x"74",x"BB",x"19",x"6A",x"00",x"62",x"26",x"D7",x"D0",x"14",x"E5",x"BE",x"53",x"CE",x"3E",x"9D",x"FC",x"EF",x"17",x"12",x"D8",x"B8",x"06",x"D4",x"A9",x"6D",x"01",x"00",x"69",x"D6",x"91",x"43",x"B0",x"71",x"9D",x"C3",x"E4",x"04",x"86",x"5C",x"60",x"8A",x"88",x"A6",x"74",x"35",x"BD",x"C0",x"3D",x"39",x"6C",x"04",x"05",x"8A",x"0A",x"9C",x"11",x"E0",x"80",x"D0",x"0D",x"A0",x"0B",x"FE",x"B9",x"41",x"76",x"1D",x"88",x"5B",x"F8",x"4C",x"FA",x"67",x"8A",x"10",x"FD",x"1D",x"A9",x"2D",x"27",x"5C",x"E1",x"0C",x"65",x"6A",x"25",x"0D",x"3B",x"CD",x"02",x"66",x"EB",x"F0",x"4C",x"C6",x"CD",x"12",x"6A",x"67",x"6B",x"C2",x"48",x"0A",x"3A",x"9C",x"C3",x"0A",x"C5",x"E1",x"54",x"12",x"B4",x"D2",x"EC",x"A8",x"B9",x"66",x"76",x"F9",x"48",x"B9",x"56",x"0B",x"43",x"04",x"41",x"05",x"9F",x"D9",x"3A",x"CC",x"F3",x"03",x"3E",x"DD",x"F8",x"B7",x"43",x"95",x"A0",x"5A",x"04",x"84",x"05",x"74",x"10",x"51",x"43",x"34",x"68",x"4A",x"37",x"25",x"0E",x"AA",x"86",x"FF",x"04",x"EC",x"56",x"44",x"A5",x"DF",x"41",x"6F",x"58",x"24",x"5E",x"0B",x"49",x"04",x"98",x"C8",x"5D",x"47",x"05",x"3E",x"4E",x"EC",x"BC",x"B8",x"45",x"2B",x"A0",x"20",x"26",x"32",x"9D",x"04",x"50",x"05",x"2A",x"E9",x"C8",x"15",x"14",x"26",x"15",x"AA",x"C5",x"0E",x"FD",x"1B",x"D3",x"61",x"A5",x"56",x"16",x"94",x"14",x"7C",x"15",x"8A",x"4D",x"0E",x"FA",x"73",x"53",x"0F",x"AD",x"0D",x"A5",x"9E",x"F3",x"7E",x"BA",x"0A",x"3E",x"4A",x"A8",x"0C",x"BB",x"60",x"B0",x"CF",x"A8",x"C4",x"20",x"C4",x"64",x"EA",x"4C",x"9B",x"5D",x"06",x"A9",x"C5",x"D0",x"FA",x"8C",x"4C",x"DF",x"1D",x"F9",x"30",x"F7",x"FB",x"81",x"85",x"78",x"EF",x"7B",x"20",x"E9",x"90",x"E7",x"5E",x"10",x"D6",x"DB",x"D3",x"53",x"47",x"2A",x"60",x"4D",x"68",x"8A",x"9F",x"2E",x"91",x"26",x"98",x"A4",x"71",x"A0",x"27",x"0D",x"A0",x"D9",x"46",x"D1",x"D1",x"0A",x"15",x"22",x"B0",x"E4",x"74",x"A2",x"B7",x"41",x"E9",x"A5",x"79",x"73",x"60",x"4C",x"CA",x"FE",x"68",x"2B",x"A4",x"DA",x"A6",x"3A",x"86",x"0A",x"84",x"9D",x"A5",x"4C",x"58",x"17",x"37",x"F5",x"0B",x"9A",x"98",x"A0",x"08",x"6D",x"DC",x"F0",x"1D",x"77",x"33",x"11",x"C9",x"99",x"67",x"0B",x"65",x"87",x"85",x"8A",x"56",x"11",x"D1",x"EB",x"44",x"0C",x"46",x"B3",x"90",x"03",x"B5",x"87",x"6A",x"66",x"5C",x"88",x"0A",x"EA",x"DB",x"10",x"B2",x"03",x"38",x"82",x"28",x"49",x"18",x"72",x"0A",x"D4",x"C8",x"65",x"0B",x"BA",x"1B",x"6C",x"05",x"A7",x"C8",x"B0",x"6E",x"8A",x"11",x"DE",x"3D",x"77",x"F4",x"4C",x"A6",x"61",x"A2",x"5A",x"DD",x"0B",x"FE",x"77",x"C7",x"1E",x"CA",x"A8",x"D8",x"A9",x"12",x"BB",x"20",x"BD",x"0C",x"77",x"AF",x"60",x"D9",x"AB",x"19",x"B8",x"26",x"A9",x"01",x"4C",x"9D",x"69",x"3F",x"99",x"9E",x"A4",x"8D",x"65",x"0B",x"0B",x"10",x"C1",x"22",x"C6",x"D9",x"28",x"44",x"91",x"D8",x"00",x"48",x"B2",x"87",x"C1",x"D8",x"D5",x"CC",x"88",x"1C",x"50",x"11",x"A5",x"B7",x"52",x"E9",x"4E",x"45",x"63",x"AA",x"B0",x"0A",x"13",x"8A",x"11",x"15",x"23",x"60",x"87",x"0D",x"AA",x"E8",x"86",x"0C",x"FD",x"A2",x"49",x"0E",x"84",x"0F",x"74",x"AF",x"E0",x"01",x"C9",x"8C",x"6E",x"C9",x"74",x"DD",x"13",x"4A",x"4C",x"85",x"01",x"8C",x"42",x"70",x"B4",x"26",x"0A",x"34",x"0E",x"42",x"0E",x"43",x"41",x"85",x"81",x"41",x"86",x"36",x"A2",x"9D",x"46",x"05",x"8E",x"04",x"66",x"2E",x"6A",x"08",x"4D",x"A6",x"72",x"D2",x"F2",x"AE",x"86",x"42",x"D0",x"62",x"70",x"84",x"12",x"DB",x"48",x"8D",x"3C",x"82",x"0B",x"88",x"5C",x"E3",x"15",x"A4",x"12",x"EE",x"08",x"6F",x"88",x"68",x"D8",x"B3",x"4C",x"EE",x"63",x"DD",x"6F",x"43",x"48",x"8A",x"4D",x"18",x"AC",x"51",x"28",x"F3",x"37",x"11",x"86",x"B9",x"13",x"84",x"53",x"5F",x"A4",x"14",x"C9",x"A3",x"49",x"13",x"98",x"05",x"AA",x"92",x"04",x"34",x"63",x"32",x"9B",x"A1",x"38",x"CE",x"2E",x"C2",x"46",x"14",x"A8",x"A8",x"6D",x"9B",x"34",x"07",x"25",x"56",x"04",x"CD",x"84",x"56",x"61",x"91",x"0C",x"CD",x"09",x"F5",x"F7",x"2A",x"9A",x"12",x"14",x"D2",x"6B",x"12",x"20",x"E6",x"63",x"A8",x"3F",x"E5",x"9E",x"26",x"51",x"D6",x"86",x"C5",x"12",x"F0",x"9D",x"F5",x"BA",x"4C",x"F1",x"A5",x"C9",x"12",x"D0",x"04",x"EF",x"D6",x"98",x"D2",x"8C",x"AA",x"44",x"21",x"42",x"26",x"79",x"D1",x"36",x"AA",x"0C",x"AA",x"F0",x"10",x"FE",x"F4",x"06",x"4E",x"6A",x"FA",x"B0",x"03",x"EE",x"FF",x"2A",x"B1",x"01",x"60",x"0E",x"19",x"51",x"F7",x"21",x"0C",x"F0",x"08",x"E7",x"F9",x"E6",x"DA",x"0D",x"E8",x"D0",x"F4",x"98",x"60",x"7F",x"D3",x"85",x"0C",x"86",x"E6",x"0D",x"4F",x"37",x"14",x"AC",x"20",x"7F",x"62",x"97",x"1C",x"06",x"49",x"E4",x"69",x"80",x"0D",x"BE",x"EC",x"E6",x"79",x"DB",x"E8",x"A5",x"0C",x"A6",x"0D",x"60",x"FD",x"31",x"38",x"0B",x"51",x"48",x"C8",x"8A",x"3C",x"71",x"B1",x"11",x"CC",x"AA",x"CA",x"98",x"49",x"FF",x"38",x"F6",x"65",x"85",x"6B",x"B0",x"A8",x"C6",x"03",x"EB",x"12",x"02",x"27",x"43",x"37",x"01",x"C8",x"89",x"32",x"60",x"B2",x"DF",x"A2",x"62",x"DD",x"B0",x"41",x"77",x"C9",x"03",x"6A",x"AB",x"10",x"E0",x"A0",x"01",x"7B",x"57",x"07",x"E8",x"D0",x"DE",x"A2",x"0E",x"10",x"86",x"DA",x"11",x"72",x"AB",x"E2",x"F3",x"6B",x"BE",x"39",x"0B",x"60",x"D7",x"86",x"EE",x"A0",x"B4",x"10",x"A6",x"11",x"F0",x"1F",x"DF",x"04",x"26",x"91",x"AA",x"B4",x"CA",x"A5",x"56",x"11",x"AC",x"90",x"08",x"85",x"05",x"5F",x"99",x"AA",x"6C",x"C9",x"8A",x"E4",x"5E",x"0E",x"06",x"0A",x"26",x"0B",x"2A",x"F9",x"B0",x"C5",x"EB",x"90",x"A8",x"E5",x"10",x"EB",x"49",x"88",x"D0",x"EE",x"85",x"F7",x"04",x"60",x"05",x"D7",x"83",x"80",x"54",x"A0",x"07",x"EA",x"45",x"69",x"6D",x"8F",x"65",x"9C",x"DF",x"20",x"36",x"63",x"EE",x"AA",x"86",x"8D",x"05",x"0B",x"66",x"07",x"A9",x"FF",x"5D",x"42",x"D0",x"0D",x"A5",x"0A",x"18",x"3E",x"4B",x"D8",x"85",x"8A",x"6D",x"2C",x"4D",x"4C",x"0B",x"CC",x"64",x"48",x"3B",x"25",x"56",x"63",x"59",x"A0",x"D9",x"A8",x"8F",x"8B",x"BC",x"C9",x"C8",x"B1",x"66",x"8D",x"90",x"1D",x"D1",x"91",x"02",x"DC",x"A3",x"DB",x"5E",x"AD",x"EE",x"8B",x"AE",x"A5",x"8C",x"79",x"60",x"20",x"D1",x"5F",x"B0",x"48",x"69",x"03",x"AA",x"FA",x"BD",x"78",x"52",x"FB",x"02",x"F0",x"3E",x"3E",x"C9",x"FF",x"90",x"20",x"4C",x"D8",x"FD",x"5D",x"A0",x"00",x"B1",x"1F",x"0A",x"55",x"D1",x"0C",x"57",x"D2",x"48",x"A7",x"20",x"B7",x"FF",x"4A",x"CF",x"1E",x"68",x"B0",x"7A",x"34",x"0E",x"5A",x"02",x"E6",x"0F",x"BD",x"0C",x"4E",x"DF",x"C6",x"0D",x"D0",x"DB",x"20",x"CC",x"FF",x"FF",x"52",x"8D",x"A7",x"7F",x"A5",x"0E",x"FB",x"A6",x"0F",x"60",x"68",x"2F",x"04",x"2C",x"4D",x"10",x"4C",x"CE",x"5D",x"7D",x"AF",x"0A",x"AD",x"79",x"85",x"D3",x"0B",x"A9",x"00",x"A8",x"A2",x"06",x"F0",x"FF",x"A8",x"62",x"FB",x"E6",x"0B",x"CA",x"DE",x"F6",x"C0",x"29",x"F0",x"F5",x"05",x"91",x"0A",x"C8",x"D0",x"F7",x"60",x"50",x"FF",x"20",x"A9",x"65",x"6F",x"88",x"84",x"AD",x"BE",x"0D",x"35",x"F8",x"9B",x"6D",x"3B",x"59",x"15",x"23",x"59",x"71",x"28",x"F3",x"DE",x"0D",x"8E",x"96",x"23",x"2F",x"91",x"F7",x"EF",x"DF",x"41",x"23",x"69",x"97",x"78",x"75",x"2B",x"30",x"71",x"2C",x"AC",x"55",x"0A",x"2F",x"82",x"8C",x"2C",x"0C",x"CA",x"08",x"0D",x"69",x"C3",x"F3",x"D3",x"74",x"A6",x"A0",x"41",x"F9",x"45",x"48",x"88",x"6A",x"87",x"93",x"A9",x"73",x"92",x"35",x"94",x"D8",x"00",x"72",x"5B",x"80",x"DE",x"15",x"AC",x"CD",x"0C",x"40",x"00",x"0B",x"9B",x"1C",x"24",x"77",x"98",x"93",x"40",x"CD",x"DC",x"AC",x"E1",x"40",x"3F",x"86",x"A9",x"14",x"66",x"A1",x"98",x"B1",x"9F",x"9F",x"70",x"95",x"6F",x"67",x"72",x"2E",x"29",x"2B",x"34",x"BE",x"C8",x"73",x"09",x"58",x"0B",x"61",x"11",x"D5",x"B4",x"58",x"A3",x"04",x"E8",x"BF",x"47",x"05",x"CE",x"42",x"4C",x"12",x"2F",x"19",x"AE",x"53",x"DF",x"62",x"61",x"4C",x"6B",x"75",x"3D",x"A9",x"88",x"8B",x"29",x"A9",x"CB",x"C6",x"91",x"95",x"58",x"53",x"09",x"39",x"D4",x"F7",x"43",x"1E",x"57",x"CD",x"B8",x"16",x"AB",x"92",x"B9",x"F9",x"42",x"16",x"84",x"23",x"76",x"A5",x"66",x"77",x"D7",x"C4",x"6E",x"8B",x"F0",x"AE",x"40",x"C2",x"E0",x"A4",x"7F",x"22",x"0C",x"13",x"6C",x"69",x"49",x"A2",x"77",x"58",x"8C",x"AE",x"64",x"2E",x"F6",x"CE",x"DE",x"88",x"14",x"A5",x"73",x"22",x"F0",x"28",x"4C",x"9C",x"03",x"7E",x"18",x"68",x"DC",x"D0",x"CA",x"00",x"74",x"0F",x"60",x"75",x"15",x"9A",x"A7",x"54",x"39",x"10",x"11",x"2F",x"45",x"18",x"EE",x"07",x"3D",x"49",x"C9",x"22",x"6F",x"3E",x"48",x"64",x"98",x"A6",x"6A",x"81",x"C4",x"80",x"57",x"D2",x"68",x"B0",x"22",x"66",x"22",x"A3",x"9D",x"88",x"DA",x"09",x"1E",x"E2",x"E8",x"52",x"90",x"DE",x"76",x"55",x"BA",x"C4",x"52",x"70",x"7B",x"E4",x"6B",x"51",x"2C",x"85",x"14",x"62",x"73",x"B2",x"2E",x"44",x"E1",x"07",x"13",x"FC",x"AE",x"24",x"D0",x"10",x"73",x"41",x"A5",x"08",x"CC",x"37",x"9C",x"0A",x"AF",x"84",x"B3",x"4D",x"0A",x"34",x"1B",x"4C",x"4D",x"EB",x"3B",x"54",x"9C",x"5B",x"58",x"86",x"4B",x"45",x"59",x"08",x"1D",x"81",x"07",x"0B",x"66",x"A7",x"B1",x"11",x"64",x"00",x"55",x"E6",x"11",x"81",x"43",x"E6",x"DD",x"2C",x"48",x"A0",x"44",x"6B",x"1F",x"C4",x"E2",x"08",x"B2",x"8A",x"90",x"90",x"82",x"18",x"04",x"1A",x"73",x"A6",x"29",x"B1",x"1E",x"B9",x"2B",x"99",x"6B",x"69",x"1A",x"D6",x"77",x"68",x"B6",x"20",x"29",x"5B",x"5D",x"B2",x"BB",x"3F",x"25",x"21",x"62",x"51",x"64",x"AC",x"6A",x"A4",x"46",x"49",x"07",x"3E",x"47",x"57",x"B2",x"E2",x"D2",x"CF",x"A0",x"53",x"79",x"73",x"71",x"16",x"AB",x"AB",x"44",x"01",x"45",x"1D",x"37",x"6C",x"89",x"5F",x"94",x"52",x"64",x"29",x"AF",x"6E",x"91",x"6B",x"13",x"DE",x"63",x"68",x"C9",x"2E",x"47",x"54",x"08",x"7D",x"91",x"11",x"EE",x"47",x"A2",x"B8",x"AA",x"56",x"1B",x"78",x"15",x"44",x"23",x"D9",x"50",x"6A",x"C9",x"69",x"51",x"19",x"3A",x"10",x"E2",x"02",x"34",x"EA",x"34",x"76",x"B6",x"E5",x"9C",x"64",x"3A",x"92",x"96",x"6D",x"91",x"E0",x"8A",x"AB",x"3D",x"6D",x"D8",x"2A",x"74",x"45",x"7C",x"6D",x"E0",x"57",x"CC",x"8F",x"61",x"41",x"91",x"1D",x"0A",x"4A",x"F3",x"0E",x"95",x"73",x"2E",x"39",x"31",x"A1",x"CC",x"45",x"78",x"AD",x"14",x"6D",x"63",x"95",x"07",x"F7",x"8A",x"2A",x"70",x"3A",x"66",x"79",x"70",x"8F",x"95",x"86",x"19",x"06",x"CE",x"39",x"84",x"65",x"8A",x"85",x"38",x"7C",x"55",x"D6",x"15",x"BE",x"23",x"E5",x"6D",x"A4",x"62",x"85",x"45",x"0F",x"13",x"DA",x"4A",x"88",x"08",x"4F",x"10",x"30",x"C2",x"28",x"49",x"D7",x"38",x"68",x"68",x"73",x"6C",x"CC",x"8B",x"29",x"B6",x"67",x"6B",x"A4",x"04",x"70",x"FA",x"33",x"A3",x"35",x"55",x"88",x"EE",x"18",x"2E",x"B4",x"E8",x"89",x"68",x"F0",x"B6",x"94",x"83",x"4A",x"1D",x"89",x"09",x"87",x"C4",x"23",x"2E",x"F2",x"D2",x"0A",x"91",x"53",x"42",x"27",x"53",x"99",x"95",x"08",x"4B",x"45",x"66",x"63",x"73",x"79",x"46",x"6E",x"32",x"AF",x"67",x"5D",x"B9",x"8A",x"29",x"42",x"A2",x"AD",x"DA",x"61",x"40",x"8E",x"57",x"6D",x"C6",x"18",x"52",x"6B",x"66",x"44",x"1E",x"A0",x"2E",x"11",x"79",x"81",x"75",x"6B",x"4E",x"51",x"26",x"62",x"39",x"AC",x"48",x"8B",x"4A",x"64",x"49",x"F9",x"20",x"62",x"90",x"AB",x"30",x"00",x"DF",x"43",x"75",x"43",x"B6",x"D9",x"BA",x"70",x"A7",x"98",x"93",x"AD",x"A4",x"6E",x"92",x"84",x"BA",x"34",x"3A",x"AB",x"7D",x"54",x"76",x"53",x"63",x"65",x"EA",x"8F",x"83",x"DA",x"52",x"2E",x"7A",x"65",x"1A",x"64",x"69",x"D9",x"77",x"49",x"24",x"8C",x"28",x"23",x"29",x"70",x"F7",x"39",x"2D",x"CA",x"35",x"15",x"0D",x"73",x"39",x"EC",x"AA",x"E9",x"52",x"4C",x"D9",x"53",x"95",x"95",x"55",x"17",x"E9",x"7E",x"A3",x"52",x"68",x"00",x"41",x"21",x"05",x"F9",x"87",x"84",x"A5",x"D9",x"38",x"CA",x"DE",x"72",x"F6",x"2D",x"6F",x"70",x"75",x"BA",x"61",x"D3",x"0F",x"67",x"57",x"12",x"09",x"C5",x"C5",x"62",x"2C",x"34",x"45",x"52",x"25",x"20",x"63",x"6F",x"BD",x"E4",x"44",x"75",x"65",x"07",x"EE",x"1F",x"CC",x"4C",x"46",x"AD",x"88",x"D5",x"56",x"45",x"5D",x"F5",x"54",x"48",x"49",x"4E",x"47",x"FE",x"6D",x"28",x"20",x"52",x"37",x"2D",x"77",x"DB",x"6B",x"94",x"B8",x"6E",x"00",x"42",x"DD",x"C3",x"43",x"48",x"7B",x"70",x"4F",x"44",x"45",x"4F",x"98",x"00",x"6D",x"65",x"E1",x"67",x"61",x"4B",x"64",x"38",x"C8",x"FD",x"BF",x"A2",x"29",x"2E",x"06",x"D9",x"4D",x"3A",x"69",x"9D",x"20",x"0C",x"78",x"87",x"51",x"5F",x"6E",x"65",x"6C",x"7A",x"AC",x"6E",x"6D",x"61",x"74",x"67",x"46",x"49",x"58",x"76",x"62",x"42",x"52",x"37",x"72",x"29",x"35",x"68",x"9B",x"13",x"4A",x"31",x"15",x"30",x"2F",x"00",x"76",x"29",x"2A",x"0B",x"32",x"53",x"52",x"D2",x"DB",x"74",x"96",x"2C",x"20",x"72",x"55",x"BB",x"1E",x"3D",x"5B",x"48",x"80",x"2F",x"08",x"20",x"25",x"17",x"25",x"3C",x"24",x"00",x"08",x"90",x"02",x"00",x"93",x"13",x"64",x"81",x"B5",x"9F",x"82",x"32",x"9C",x"34",x"23",x"4F",x"28",x"AD",x"29",x"EA",x"68",x"50",x"59",x"CA",x"8D",x"47",x"48",x"EE",x"74",x"47",x"31",x"37",x"EC",x"AD",x"30",x"2D",x"32",x"68",x"50",x"25",x"55",x"B5",x"47",x"B2",x"20",x"93",x"57",x"94",x"2D",x"C2",x"F5",x"49",x"50",x"48",x"8B",x"4E",x"3A",x"7B",x"43",x"CA",x"65",x"00",x"23",x"A9",x"2A",x"4A",x"71",x"97",x"5C",x"16",x"48",x"41",x"D3",x"53",x"62",x"7F",x"43",x"55",x"D0",x"C7",x"45",x"44",x"43",x"FE",x"7E",x"25",x"52",x"9F",x"F9",x"03",x"3C",x"20",x"80",x"00",x"58",x"93",x"49",x"4B",x"7C",x"4F",x"CB",x"72",x"CF",x"25",x"73",x"65",x"FE",x"46",x"6F",x"75",x"6E",x"BD",x"CB",x"66",x"69",x"5D",x"EB",x"3A",x"20",x"06",x"18",x"2E",x"A1",x"80",x"3F",x"FD",x"1C",x"6E",x"81",x"FD",x"0F",x"80",x"81",x"AF",x"DA",x"D6",x"D1",x"03",x"49",x"50",x"52",x"17",x"2C",x"55",x"2E",x"DF",x"4E",x"59",x"0D",x"6E",x"3D",x"A7",x"06",x"B0",x"05",x"22",x"2B",x"4D",x"51",x"52",x"4D",x"41",x"77",x"20",x"55",x"E9",x"29",x"4C",x"34",x"EF",x"59",x"00",x"3D",x"D6",x"54",x"12",x"A5",x"88",x"E8",x"70",x"B2",x"65",x"64",x"D0",x"3D",x"A1",x"80",x"20",x"4B",x"42",x"E2",x"2F",x"39",x"00",x"56",x"E4",x"8A",x"6F",x"4E",x"79",x"09",x"31",x"66",x"1A",x"43",x"39",x"78",x"10",x"4D",x"BA",x"78",x"69",x"8E",x"75",x"6D",x"76",x"72",x"5A",x"45",x"64",x"61",x"62",x"6C",x"1F",x"5A",x"65",x"63",x"74",x"EB",x"18",x"C2",x"73",x"F4",x"00",x"57",x"D9",x"FB",x"95",x"2F",x"2A",x"65",x"85",x"6F",x"A2",x"72",x"40",x"A3",x"20",x"01",x"24",x"8E",x"47",x"55",x"A3",x"4D",x"69",x"C0",x"42",x"45",x"53",x"89",x"43",x"41",x"52",x"BD",x"20",x"46",x"4F",x"55",x"56",x"7A",x"2E",x"00",x"DF",x"30",x"31",x"32",x"33",x"9F",x"F7",x"36",x"37",x"38",x"39",x"C1",x"C2",x"C3",x"FE",x"C4",x"C5",x"C6",x"2D",x"32",x"31",x"7F",x"37",x"E8",x"33",x"B0",x"36",x"34",x"38",x"E3",x"C7",x"0C",x"09",x"0A",x"10",x"40",x"F9",x"50",x"A0",x"D0",x"3F",x"64",x"A6",x"52",x"87",x"0A",x"00",x"33",x"4C",x"0C",x"40",x"12",x"44",x"14",x"1A",x"70",x"11",x"01",x"7C",x"A8",x"00",x"60",x"0E",x"03",x"91",x"68",x"02",x"8B",x"86",x"66",x"09",x"4E",x"62",x"40",x"F4",x"55",x"25",x"06",x"38",x"22",x"0E",x"A2",x"01",x"C3",x"02",x"86",x"03",x"56",x"01",x"05",x"D2",x"2D",x"17",x"B0",x"08",x"07",x"09",x"E8",x"04",x"14",x"47",x"15",x"06",x"16",x"17",x"AF",x"18",x"35",x"19",x"74",x"1A",x"03",x"1B",x"7A",x"1C",x"0B",x"1D",x"06",x"F4",x"1E",x"1F",x"A7",x"0D",x"20",x"21",x"D7",x"22",x"07",x"27",x"E8",x"01",x"31",x"03",x"32",x"0E",x"33",x"7F",x"34",x"08",x"3C",x"06",x"F4",x"3D",x"3E",x"AB",x"01",x"3F",x"09",x"40",x"3F",x"41",x"0E",x"42",x"07",x"43",x"FD",x"46",x"06",x"47",x"E9",x"48",x"AD",x"08",x"49",x"03",x"4A",x"04",x"4B",x"FF",x"07",x"B0",x"4E",x"0B",x"8B",x"14",x"42",x"49",x"47",x"53",x"54",x"3F",x"4D",x"4D",x"30",x"16",x"FF",x"2C",x"B4",x"BB",x"EB",x"58",x"90",x"F9",x"56",x"72",x"31",x"C5",x"15",x"D1",x"13",x"F1",x"46",x"C6",x"19",x"89",x"E8",x"0F",x"E1",x"76",x"48",x"87",x"02",x"8C",x"96",x"43",x"06",x"04",x"1C",x"F0",x"26",x"29",x"6D",x"66",x"62",x"61",x"4D",x"7F",x"45",x"47",x"AD",x"51",x"2E",x"A9",x"26",x"46",x"41",x"54",x"33",x"32",x"F9",x"C0",x"20",x"0E",x"1F",x"BE",x"77",x"7C",x"AC",x"FE",x"22",x"C0",x"17",x"78",x"56",x"B4",x"0E",x"BB",x"07",x"00",x"3F",x"10",x"5E",x"EB",x"F0",x"32",x"D6",x"E4",x"16",x"A3",x"CD",x"19",x"EB",x"FE",x"AF",x"B2",x"E2",x"48",x"59",x"35",x"50",x"68",x"42",x"28",x"4F",x"A8",x"A2",x"56",x"A5",x"D6",x"2E",x"82",x"31",x"EE",x"0D",x"3F",x"4E",x"ED",x"4F",x"0F",x"47",x"53",x"F2",x"34",x"79",x"21",x"11",x"5B",x"63",x"65",x"5D",x"F3",x"32",x"AC",x"2C",x"36",x"EB",x"61",x"2C",x"38",x"35",x"31",x"E4",x"30",x"9F",x"50",x"2E",x"43",x"96",x"05",x"53",x"6A",x"0C",x"20",x"34",x"59",x"4F",x"28",x"8B",x"6E",x"CB",x"58",x"26",x"54",x"4B",x"55",x"35",x"D2",x"D4",x"A8",x"12",x"4C",x"D2",x"43",x"4F",x"4D",x"50",x"F5",x"55",x"9B",x"45",x"B2",x"8E",x"4E",x"44",x"3D",x"54",x"52",x"59",x"20",x"7D",x"94",x"49",x"B8",x"4E",x"5B",x"50",x"52",x"45",x"41",x"EB",x"44",x"59",x"2E",x"0D",x"0A",x"00",x"FF",x"61",x"A0",x"01",x"F8",x"99",x"EE",x"0F",x"08",x"3E",x"14",x"85",x"53",x"AE",x"93",x"4A",x"F9",x"C2",x"38",x"02",x"0C",x"38",x"C0",x"23",x"12",x"46",x"44",x"C5",x"49",x"5B",x"4B",x"4D",x"45",x"47",x"41",x"36",x"35",x"FF",x"59",x"53",x"68",x"30",x"D0",x"80",x"50",x"08",x"BA",x"32",x"69",x"74",x"0B",x"7A",x"26",x"22",x"28",x"62",x"63",x"6C",x"64",x"20",x"1B",x"D2",x"CC",x"55",x"D7",x"B4",x"65",x"06",x"8E",x"36",x"29",x"1B",x"4D",x"D9",x"34",x"DA",x"05",x"A8",x"64",x"EC",x"45",x"26",x"AE",x"09",x"63",x"85",x"04",x"4A",x"54",x"00",x"65",x"09",x"D5",x"D3",x"58",x"52",x"04",x"03",x"02",x"07",x"F5",x"06",x"08",x"9D",x"75",x"4F",x"51",x"08",x"83",x"84",x"02",x"01",x"0D",x"30",x"18",x"5C",x"34",x"0D",x"37",x"BD",x"B9",x"9A",x"A2",x"64",x"16",x"65",x"56",x"7A",x"6B",x"2A",x"8E",x"6C",x"BD",x"75",x"C8",x"88",x"B9",x"1A",x"8D",x"74",x"D9",x"8C",x"77",x"D2",x"79",x"20",x"43",x"D1",x"CD",x"D0",x"E8",x"60",x"01",x"3D",x"02",x"E8",x"A1",x"00",x"03",x"85",x"30",x"31",x"6C",x"06",x"28",x"00",x"A0",x"C0",x"02",x"F0",x"07",x"A9",x"E6",x"BF",x"92",x"4C",x"56",x"6E",x"60",x"A2",x"19",x"B5",x"02",x"9D",x"FD",x"95",x"79",x"CA",x"10",x"F8",x"BF",x"00",x"A2",x"D0",x"85",x"F5",x"02",x"86",x"03",x"6F",x"0E",x"5A",x"D2",x"41",x"AF",x"96",x"04",x"B0",x"DC",x"AE",x"79",x"A9",x"05",x"A2",x"03",x"A0",x"BF",x"20",x"BA",x"B4",x"4C",x"C0",x"FF",x"D5",x"F4",x"79",x"49",x"44",x"22",x"D8",x"99",x"15",x"D1",x"D0",x"88",x"88",x"36",x"AF",x"66",x"22",x"DC",x"59",x"11",x"D1",x"00",x"C0",x"90",x"D1",x"CC",x"88",x"88",x"44",x"B9",x"30",x"3B",x"99",x"E6",x"07",x"88",x"D0",x"F7",x"18",x"AA",x"98",x"29",x"0F",x"99",x"68",x"03",x"F0",x"0C",x"8A",x"79",x"67",x"03",x"99",x"68",x"03",x"A5",x"9F",x"79",x"9B",x"03",x"99",x"9C",x"03",x"A9",x"01",x"85",x"9F",x"A9",x"78",x"20",x"00",x"01",x"4A",x"AA",x"F0",x"09",x"08",x"06",x"9F",x"38",x"6A",x"CA",x"D0",x"F9",x"28",x"6A",x"99",x"34",x"03",x"30",x"05",x"A5",x"9F",x"86",x"9F",x"24",x"8A",x"C8",x"C0",x"34",x"D0",x"C1",x"A0",x"E7",x"8A",x"4C",x"9C",x"01",x"40",x"00",x"79",x"69",x"80",x"0A",x"10",x"0F",x"06",x"FD",x"D0",x"08",x"48",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"68",x"2A",x"30",x"F1",x"70",x"01",x"60",x"38",x"85",x"A7",x"AD",x"29",x"01",x"D0",x"06",x"CE",x"2A",x"01",x"8E",x"E7",x"DB",x"CE",x"29",x"01",x"AD",x"3A",x"3A",x"60",x"20",x"1A",x"01",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"66",x"A8",x"CA",x"06",x"FD",x"D0",x"06",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"E8",x"90",x"F3",x"F0",x"E1",x"E0",x"11",x"B0",x"51",x"BD",x"33",x"03",x"20",x"00",x"01",x"7D",x"67",x"03",x"85",x"9E",x"AA",x"24",x"A8",x"10",x"09",x"70",x"07",x"A9",x"00",x"20",x"05",x"01",x"D0",x"25",x"A9",x"F1",x"E0",x"03",x"B0",x"03",x"BD",x"A2",x"01",x"B8",x"20",x"05",x"01",x"18",x"AA",x"BD",x"34",x"03",x"20",x"00",x"01",x"7D",x"68",x"03",x"85",x"AE",x"A5",x"A7",x"7D",x"9C",x"03",x"65",x"FF",x"85",x"AF",x"A6",x"9E",x"B1",x"AE",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"CA",x"D0",x"F1",x"86",x"A7",x"F0",x"99",x"4C",x"0D",x"08",x"CC",x"F2",x"01",x"00",x"0B",x"08",x"13",x"02",x"9E",x"32",x"FC",x"30",x"36",x"31",x"07",x"00",x"A5",x"B6",x"8D",x"53",x"D9",x"29",x"F8",x"09",x"06",x"85",x"01",x"BA",x"FE",x"8E",x"A9",x"26",x"BB",x"79",x"2D",x"E4",x"6C",x"5D",x"58",x"47",x"48",x"F7",x"62",x"A2",x"DD",x"19",x"BD",x"47",x"79",x"95",x"02",x"CA",x"10",x"F8",x"68",x"50",x"52",x"4F",x"50",x"2E",x"4D",x"36",x"35",x"55",x"2E",x"4E",x"41",x"4D",x"45",x"3D",x"53",x"44",x"43",x"41",x"52",x"44",x"20",x"46",x"44",x"49",x"53",x"4B",x"2B",x"46",x"4F",x"52",x"4D",x"41",x"54",x"20",x"55",x"54",x"49",x"4C",x"49",x"54",x"59",x"4D",x"36",x"35",x"55",x"4B",x"45",x"59",x"42",x"4F",x"41",x"52",x"44",x"20",x"54",x"45",x"53",x"54",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"EF",x"01",x"0D",x"08",x"13",x"57",x"2E",x"59",x"01",x"08",x"0B",x"08",x"37",x"01",x"9E",x"32",x"30",x"36",x"31",x"00",x"00",x"00",x"BA",x"BD",x"F4",x"08",x"9D",x"FC",x"00",x"CA",x"D0",x"F7",x"A0",x"35",x"4C",x"A6",x"08",x"4F",x"BD",x"5A",x"08",x"FD",x"9D",x"48",x"07",x"CA",x"10",x"F7",x"A9",x"FF",x"FF",x"15",x"5B",x"8D",x"16",x"D6",x"4C",x"57",x"08",x"7F",x"06",x"3A",x"55",x"37",x"13",x"D2",x"C7",x"C3",x"9C",x"0B",x"0E",x"64",x"BF",x"CD",x"0B",x"C8",x"5E",x"0F",x"15",x"ED",x"05",x"03",x"E6",x"0C",x"19",x"2C",x"1D",x"75",x"38",x"F0",x"0E",x"04",x"9D",x"17",x"42",x"1E",x"AA",x"01",x"2A",x"FB",x"0F",x"8A",x"0C",x"B5",x"07",x"AB",x"8E",x"57",x"15",x"10",x"EB",x"12",x"13",x"08",x"09",x"06",x"14",x"7E",x"20",x"AC",x"52",x"4F",x"50",x"F5",x"96",x"36",x"35",x"55",x"2E",x"4E",x"FB",x"5B",x"4D",x"3D",x"4B",x"EB",x"59",x"42",x"DD",x"4F",x"41",x"52",x"44",x"20",x"BF",x"45",x"53",x"54",x"00",x"DE",x"04",x"04",x"08",x"00",x"0C",x"80",x"C0",x"00",x"00",x"84",x"D0",x"40",x"00",x"48",x"80",x"04",x"40",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"B9",x"9C",x"09",x"99",x"E6",x"07",x"88",x"D0",x"F7",x"18",x"AA",x"98",x"29",x"0F",x"99",x"68",x"03",x"F0",x"0C",x"8A",x"79",x"67",x"03",x"99",x"68",x"03",x"A5",x"9F",x"79",x"9B",x"03",x"99",x"9C",x"03",x"A9",x"01",x"85",x"9F",x"A9",x"78",x"20",x"00",x"01",x"4A",x"AA",x"F0",x"09",x"08",x"06",x"9F",x"38",x"6A",x"CA",x"D0",x"F9",x"28",x"6A",x"99",x"34",x"03",x"30",x"05",x"A5",x"9F",x"86",x"9F",x"24",x"8A",x"C8",x"C0",x"34",x"D0",x"C1",x"A0",x"C6",x"8A",x"4C",x"9C",x"01",x"04",x"00",x"08",x"69",x"80",x"0A",x"10",x"0F",x"06",x"FD",x"D0",x"08",x"48",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"68",x"2A",x"30",x"F1",x"70",x"01",x"60",x"38",x"85",x"A7",x"AD",x"29",x"01",x"D0",x"06",x"CE",x"2A",x"01",x"8E",x"E7",x"DB",x"CE",x"29",x"01",x"AD",x"A6",x"08",x"60",x"20",x"1A",x"01",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"66",x"A8",x"CA",x"06",x"FD",x"D0",x"06",x"20",x"1A",x"01",x"2A",x"85",x"FD",x"E8",x"90",x"F3",x"F0",x"E1",x"E0",x"11",x"B0",x"51",x"BD",x"33",x"03",x"20",x"00",x"01",x"7D",x"67",x"03",x"85",x"9E",x"AA",x"24",x"A8",x"10",x"09",x"70",x"07",x"A9",x"00",x"20",x"05",x"01",x"D0",x"25",x"A9",x"F1",x"E0",x"03",x"B0",x"03",x"BD",x"A2",x"01",x"B8",x"20",x"05",x"01",x"18",x"AA",x"BD",x"34",x"03",x"20",x"00",x"01",x"7D",x"68",x"03",x"85",x"AE",x"A5",x"A7",x"7D",x"9C",x"03",x"65",x"FF",x"85",x"AF",x"A6",x"9E",x"B1",x"AE",x"91",x"FE",x"98",x"D0",x"04",x"C6",x"FF",x"C6",x"AF",x"88",x"CA",x"D0",x"F1",x"86",x"A7",x"F0",x"99",x"4C",x"0E",x"08",x"CC",x"F2",x"01",x"00",x"0B",x"08",x"FC",x"9E",x"B2",x"30",x"36",x"32",x"FE",x"0B",x"78",x"47",x"77",x"53",x"84",x"2F",x"BB",x"63",x"41",x"85",x"47",x"A9",x"7B",x"F5",x"8B",x"21",x"D0",x"8D",x"9C",x"D7",x"FA",x"07",x"5B",x"20",x"93",x"22",x"04",x"5A",x"0A",x"81",x"FF",x"BC",x"E8",x"A5",x"03",x"01",x"43",x"54",x"0E",x"00",x"A2",x"50",x"52",x"4F",x"50",x"2E",x"4D",x"36",x"35",x"55",x"2E",x"4E",x"41",x"4D",x"45",x"3D",x"4B",x"45",x"59",x"42",x"4F",x"41",x"52",x"44",x"20",x"54",x"45",x"53",x"54",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00",x"00");

begin  -- behavioural

  process(clka)
  begin

    --report "COLOURRAM: A Reading from $" & to_hstring(unsigned(addra))
    --  & " = $" & to_hstring(ram(to_integer(unsigned(addra))));
    if(rising_edge(Clka)) then 
--      if ena='1' then
        if(wea="1") then
          ram(to_integer(unsigned(addra(14 downto 0)))) := dina;
          report "COLOURRAM: A writing to $" & to_hstring(unsigned(addra))
            & " = $" & to_hstring(dina);
            douta <= dina;
          else
            douta <= ram(to_integer(unsigned(addra(14 downto 0))));            
        end if;
--      end if;
    end if;
  end process;

  process (clkb)
  begin
    if(rising_edge(Clkb)) then 
      if(web="1") then
--        ram(to_integer(unsigned(addrb))) <= dinb;
      end if;
      doutb <= ram(to_integer(unsigned(addrb(14 downto 0))));
    end if;
  end process;

end behavioural;
